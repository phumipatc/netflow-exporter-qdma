`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
dXrgiZCp8UsbYFNAQXZepTXFlYCtZOjh260C3fwE2kGd7eQu0YYlfnHl84NGhOAPkKv72LfiQrp1
D0bBr/gB+ghb7QJsO2a5wqDkKGC56TloCpOrIKF3bMp54e+N9wxxOcX4oxNTWWwZONV9xjs18utc
fIdkxzPuQxgJsZQ4gKOtFlgktfcYHSFysXWp1HIxeOln11Txh/t/4ykGEdk47k8EisPMyDQJQ4mR
54lojqD10DzEU2efKXyR8ffTCK8pW9Td7yodhJzYzvdaDz7ul1D2JcsJBp1/8CrbDjIX2CkEOFpq
oXP3yNuZXVZNr95pKtZ7a6XlmR47jTTYdcxgwA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
GuS7S54ZrAFeN2mdDVw4MZfvc0Sx4qrjbbtmn3qA77xwH3rJ5uvRPQWS9Qt9kwBuPxBPARFYKdY3
fcsHTywdJIa5Y0tbPakTpoQQyT8OwQcj1Tp3plPwqEWbSiWsf4UQGe6dRTgF4UfWRtYwaq7wIKsm
gCVxRFOcNvkynr061kE72ZFakopSBQSaJtTNJpBmB5HjMDcxgae3cyTrukH1+U58NoR3XDkwyypM
YDzonO+xUfAUfdDR7z3fUPlCr7ubvsWwki+ndNJarGcUewkXyI1M8ZYve14CEeHRAmmtflRJIzMQ
PH1lY1zqpQbnz0UxYp8KW1zYB6Lrf2Y5dR90VAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
SctbpSY0YT7+L711CObLnbmp/N5a/DzGwssFc+ZKj+JQwFYTh4hmPgzpQYgdvBeBOe4nrhJVKhE/
OOHO5W+xow==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
IT6ZiNUm5BF1bQuQ3SB+Fm+ZMzrCmLfmUNzGmPQ6Ge1k2vp9H2b9HF5MwxCElPehfatPQO9PsV2U
XGASNRYQolKE3z+EvzLAYVpkZWYF5pY6JhJzO0cU7l1pay3x0ehXIQt3Q0hQvS8Pg/7GTzn3oBe5
iRU8V/CZgczdM9MYKTo7vu/rBRRvJWPyheLQ+eTGyoL08vrUi5xUhxFK3v3NUhXQFtk9pzre8QRv
cX7hwwMjQO2MH025wTbI3P4dHQC3N+VNeN8knxtgfB+8a7H6DL3JRi9RPGCSW/peX5VOKjysJvTO
FWLl19/tCEE2rV17tS5gf7BczqJo8LR39kds5g==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
P0ehh15jAdAXY6IUWlEQlsdKlefuYn+9qUV7zNO4i+P9UOPfrdt7/7E0ZsSDaLKSPxztNjtUqiX3
WIlhZdkpN/UklalkejsxwK24VSw8g/ofeuDDxRR1FyLvu+oe2BqjsPObBFjivPFBlt8c5rgrLPWf
g6W9eZdx6LG8J5JYZXfx/alzegazclci1lMXmLuKiHsPf/FDRmHmPAnAudJkfHryTHNlRNnuJUk7
rTHmVa700pAn9aUVuo8kZ8+yxoqYmbwjgfDuabViqwpohPhErXdcpa56nl5/09qHNI1zB+jO1zs1
dK0+asQB15sByRV+I5f6UtUlugpH1lxStxAQCg==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mIQUoljSgJbaO9nDzmkfw/axQzhzo63ekQwezHbMIA+gf6NX5f0uf2xRueyuQgYbOYp4v+/L7+GC
fjEthCumqOhDkmDW7IKhqKhf4ZRmiC7+WljbPyf/FHgtkKAjsmYWEiQDWp59/jY+smzigSeGFUYf
Vu96zLNxJ3pjbKiOABY=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
G2KTZ93n+PxAfw2zfnA1COabZno1DRWn0WErnZMXT9uCatPRkkfxbLXrLwOELRAZVLsDiWR2713W
nmUyqfMQWMnSjtML6cbSydef2ppz9fN6DwIGMufcuypUdy6OrAFTeIt7LkrPpVC7aqWgvMOKZLQK
qu/ILtLzYwfEAtl5hX5/e0I/ADjPah5TKxSzFk6Q3Rddqp2qcTc2zkrnpA+0DiqK+/r0qWH0IMbn
Vn07LiixWV5OyfWrSLHMmsx2gwR728MKiwkZCD3Rt65/fl1mXfQm+q2tr+eaDxmU0fzvFaK6ct2y
46tpqf8vOlSJ0klBX1VsoHtgGcP0HELExsjKFw==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ihF7THQrde8/5fKBj4PNaAyrdLLezirPwjVM0qEROgu8Xewo//jwFzLP5WaSOkI+ZHFjmejkkOWB
3xyxiEIZ2+bvMCjklc1mGbxleYJ/zUr0Wn7SrwtNIK5GtrtR3u2z0wWYSQxmMguJZSWZSkUJKr2q
hwDrfvu36x0M2vBOD/KHEVX+htbbDDBGjYWFXlAFl0xymU8yZZIVYfTiCUqqIy6E5toDg7Ws+5S1
6E6VCv5J+aIpt9hwe5kmHnvkXcamG96Sg23XlVPCr20M3Z+VUTsTgJGZn7PgYsKv6D1mqzoVBrSx
Prj6O/LvBjASIBE49zTRE/G1cPNUVdWiqEgFsw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
B7ExKxhazC7ZPZBruibWY//nhQ3KB7LnX/NjjNuvPu8X7fffms/t/Qpwx4fQhrHXoN+MUeduogqe
7ji3bpTW+yiB804QRzrZuvoxTbRedxcZcexDC4kuLvaRI5WRhQYlaix6vp9v0TNUP6VLAWTcxS1B
jK/PEXCKHXZylKGig6g=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
R72hR7jVo3GwTawy14vLHQzaJqWicpvVYav3UoTxx3iQC6YkH2sOwCG0JySKUypzQj5+TRSXC+sL
UII0q/KlKzhdq8/8/0bEGKX5kX1aoZU78SRHaB2MhUpO7jXIo2VwWTss9gKEKdiPvrcVOBg0wY7/
1N4wPHKnJITxOp3IqeEdc8ZXFZFKFaAhGa32cEoDZ+F9yfUpP+2RbWTp+HvlJgoB8TpE2Gt0wjWG
rHIJXA2Cz/l2gJyRwTU53nrZFwB7LCTwc3s333dM8PTkI+7mv7mhMTDT2SW79eyGpSkXUznJI6j2
eRI+jZF9Q6oakV8mIQoxwfMQy12RN8Vi+zX1ag==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 31264)
`pragma protect data_block
yadlYB4YI477RiEZPtEHoeWlCoXQxWwf7aQSWgIy+670ontQIC4YENgePyaYfPNGAWoVzHFX3w3X
VjZtpH9dv3/ISlgiYsXp00SnvY+B3UQAjKdAsD5o2XsL3G6aE0nMLjqsbklDXLs7zq6EicD+3SPf
L0AUMSF1DUKKh4gMUBxIxIr7GvD4pyoa7cEmA0X1DrogsK7BnyKZamOYM4PwyCE5mxMQaHl5y6Fb
bOo1ouTgsYkBK01UCNe3X7BFqpD9fjyTOLSmyMoObh/gdSN5o3NbVkvpr6ZFuPe3l7/bFLArCk9o
F48/86HRiHxKGFRR3tpye9PvQp97dz6JzgkGxP8w8Sn4Z9lf9Og0q1JvFC3OjSMRD1yXV1E4ARL2
/nSRhncQA5EGS2V8v0H2BXRZFsl2QIjNcPxRcHud+hlplbIllmxtJn1OiYZ9rj+2T5jFXybwkCf8
91RYeCqg+aZ4dqfuKaRS6BU6D1WMLYpIgnqYwamAi7rLQVBpjRWZseYAULDUyZXiat4SBQCNyBRP
7Mc8uH3ztjQNiYFpO9Psto2rA3X91MDpYCl4yNmfe4NPww2JRnakKXDW2GyeixOHW3gLdjTwEkPV
0YcK9vOMqmuqfvTyeYfzo/7n47yQrDTopVRQ34kV9NxcgKs+8mCChLc8V48FLiXqvulbL0ZiW+Tc
s6A/XVaM8gDBuIeg54Hs7NlEUJEnb6fcmjmu1hxanpBAD5mJMkAvilIF5DqrDoLxJy196Lpy34AY
2mRvJ/cbHD2M89Bm5iHYsRG8eohaP2Z5krqMQ5MisxR5HHupVitszGVXl2u3OPl+SgqTKvFyoEFA
SNAtjOZMBACgExURMo1ko7Qq/x/lhUNHSrYIaZooNWE9GluhEkEopfzuOUh8qZ2OJwKpHe1zlz+Z
fygFlGbgd+TO+pdO7XcAfdCHW8sGlqehgamR63kTC7thmAqKR8G+dKl/7w3W6cncdcMfdVGY7glT
VYLEHMdO67SiREAThlASs+wMTdiBZtrQxxF216UNoH+VEtSh5t9y6O9gYxXgrML7PBbN1B4JX1Hk
vnmu0i8gB827hfJlE1T8lk0DigmYtOzTj4y/Dv6RA9ksGPoJr8uHBLT9lJ+NxzQkFkaDX3qBhbQC
TT3culuwbV3dREyvcTQW0EzOPM2ldxON5msn8TjAPu1ntiF4fvFg7s3nxwXTMOUC98+O1ggCAGgB
n4mXV11QhLsKktov5dH/LNtvZFyCppUz3Qn/ewzg6B+j7j4xR2un/lNcNoY2bI/AjaDkU6inSVN3
39tluXj9lPf35Vx4De5XdGmJJTC6wubAdty0ZxZJKPulamFNYZ501iTrXrk7+MrfP9Z3fHj1zyKD
lDqtxKVvdoxw4Jey8LvXVKBqRmUb9U1P7Z53EaMMOvG44Gf3OK+wYC1qV0vk2dtbTjaXvMYrYMU0
VsR3/JOWkhJKb+7KGIagOHUTx4vedHR74YAkkABuig9awt30JuLKZKvuTpDJ1/k/kjn5JMpZFJhU
bzs+In4sORzaQi1TtZD9JjZm6/Tz3dKv3I7nj9Peza+kAVoZIaXrlgqlyJLPuvztRydqsLLPm3f3
ghs7MUUVv/aq3Zie4XHTf+aMHfAhWv4/0OUWZ7lo+PSDntlofU6nmXLMGNnIQzAM9pG7Tzh9i5RP
A0DNbijaEWxQMxMl8leIPJoNTPSyRiT1ct7E/Y2Tz8zKvm2jXpTB/jYxrnoHVNiyhcJNlOQ5ZtvK
xgrQl4gxg8RgzzTijCbg9h/B8jpEkTJR3KWbvuBZ4gL4etea8B9Ao3GV1n/CCzhvEdJJgY+QtTWV
b1v03yZF0Q6H693heocM8h5Og6cQ54b+j5YUSs4w4Vb5CO9/qlupzw28i9d38bBZ9+O3RNlK72VA
iqULuJXBglxjcoWoYAhrT+Swo7jtQi4tuP2bpDqlQlo2vN8BDBXL9AV8VlhpF1GrjxP5cwQ6X64a
nfevGf+bZjRvci3P/wEO+qWzpG8eYjaGtcC84omDkfN9UHfol4ehvaLZeeQN3Bt43Kftud7vBF7q
ugyv5fFs4vSJiMCFkTiXbXlCBgHe2clxrXJDVt2KXdifpvJOMHoUI8STE8U2p6GlmUrqGe1UabTH
8SsYPTPZtu3Xwhwnvg6mJOtYmye+PNlDcO1o9WjlkWnea6BTcLP5WB0J9NSNDDg97JrTASJ2KSLM
VsK+yDKwwXbgcgP/awkhb8iyGIt7fA+MnHvFkPgfYsJmcPx4mysRntP9JtHxdFF35/d5aqrFkl3i
ssyKig0uOyq+VR1hhp5pckzFiCnpfLsayA+h/uoetmujLe4u7kQSADObG61LcZhEtd4dcFlUqVpT
eE953xkjKmabcYBAaAOcqZtkfjiEuTBL/KlCsz2R4Gh8hsT0xKgRgJbYwKn4aGp3b0EygWr1XMNr
VXM1WL15/igKChBOiz+/2CAQbSEa1BeLPT7DvG0E25KYFbmzH5QeoI0cx4qKYrKbTKwQVGdhnZQA
NSoz2qK9VP23N/eHwCLH7Y600EVETUH1pDrngbAD74HOqNn+wsjTzvPojkUmpRsu5e1ofCplm9K9
Qa+fbH8k+GuiSwfcDAMXrmbl0ixEJFinvG7+q9vZJw3d3ygXL7K7H5dGon2HSw+WzXKpNaqZPr04
wZ7BmK2kUjpXxvuNZvXUVF0T5Ro+JUF+66rOqKbN26885NNP0F0gP+WbqrWt8fXDF2baHSoX9zYQ
Yr9HMzI+naoA9BNbl0wiSwv7Y8/ljjg+u/QJ4HTdkEai9U+P8WXTDm0+ApujEtduCdaxwruEMrqP
x33xjd1+ZFVRAZdVyC+oAUIbALHCTgOaakCTbUn369ikWzyVutTGd9zXGuAehw5UlzG51Ug21AQ0
VG5kOHplV+2U1UOKeJbPp6u3/paryXmBYNiCExvhXT5MA5350G6wDiAyrPgM7/XY9Iwxj4OtiNC5
selPnhXIbLtczKa90R0/32NDOJxz11ImaZwdg7XecLHkasjSJhdjeSRvqDQ9jaZj3EdEPg4auuMX
Gd1QuG2oOLbChx9/nuxQHS4sMC3Kht2sqpICIWKTW/l725KqNDkSDkRPqlGI0lbfL6/+oTJ3idfh
Dd03YWfJpq4KPGXoa/dWlq5YdpPxEcCsYv0ETgAKV6TS0SxiJUBDQPZoWavrjyNpwjRCdxtGsWFM
FEMcpgC4SGoOHTr/7Fi9G/dBlmRsdwI0ikZ4a0jCnu6w76J1kPl34LAV3fqsaI9Cu28CCP79iqKW
2a+S8wLQBQ9hItJH3mlJVdrShO9RJpleWzwz77wVzHoNSQnjJEX0UJLTIo2IktG8kq8nVyGDYVQD
ydIH+RVd7MwAbGHKhYfe/7kQ5RbdXKuQHZjHwTA+lXU2Ql/OAvEpT4IHnohrBzEUbG9YlBr6Ed/u
5XfNTgDAtBPh6+OtOXOMDGk45bnZkjlqDBO47LaKq9KfLo9mnvz0rrqpzDsXo+nPKVo5N79aatZO
2JGc/hOBrqrzmChuJGvkepetVnoLfMHn5n/jHDjgk9hQYNPGRxAibLPwUyiDXbrCPD2T41gikOf4
WT82e41aUY1MsevZQpPP/3UyHZ5sCNP7tLPS0gknD8taLxvsxAH5fRvwC5D+cTZGU5svVTlTGIGy
f95z2kbB5O1wjIBV5dNH1iwhGmL5SZii8YqTYeEPbRy2rJR0OQqHbENTwVF/0gbnfKIDsPIFJXbc
7nR7XwaSKbD5mZ4IzBCXajG2W34IV/XzBKNM/UUC8kQrF7vAwec2/183KuP/C62wO93+0ooTDq9L
O764npFPbWt8DQ2mQa5WHoKladga9KIZCNB5jHZnV1AJbHu/+AWW+ZaIzXrBrbrKaTMfJN5gKraF
mQqaVvEjP6w0FnwU7dS2i2tYhOzQrA9hnePq7LaIkBMzrifEW/D1yIv97B00P0RQFfb4Bo6kh59+
1FdkBjX5Mr2bFpvH/8HRgKIzmrCUEgPREdGQbSuCHtnLKhCd+m74g2os59OfXFe1TE3JOjXIqiU3
sAl2DLQMYdrL2Eku3Hlvoxs6Ody3uXGH5XRxS49ee76Fy1DzRiZPTELcCcI+WnfltmElnVYArtJQ
Ga2GBXW6GH3541s+Q3fq/hMDDyn477J1ERlwe153X8jNmfNoRC1MF5kfh3SoOuOue+r/fwmVD3bD
DImBTmwioqoyy6IMJ9g5aSis+xhjN88MCcZ32tm4A3FMjey/0Db0gRnzcfZYHR5IwwgwnP6Ie7Bm
scC+MYhD1cWoYVZBg2/oVWqhhi7dzA5LiqyPMHhSp9pWfucPGpuJmGFfLHP/qQxC/eQMcacjMyu1
gHHp0tvBfpnSLkj4X6ld5vfvCeDcTMVyOHlKHDs1fC/epzGDYP095PVguYw1bbSMdq4h/mCYjU+6
AX5T4ckwyCEt1qh1+YbF/9DNVHBN3jhvT2OD+75znS8R5/HZIEWVBsJye47TbhizuN/BP8Og0d5m
w6J1lnhd/Xy+Z8UkcF0BHJ/PuYzJGHqGNtKed5icLMowf0F1TCbq/8Ymuw73CYVgUvh3LCwa/tQH
GvlIWb5C28ivzYr4ua6eeLs4gu9EM7qKMXr/pdZ6c+0mUXR4cKlYF8HkyL76l5ASe9P/qM853HXf
OToIYKeub/cIlwN/Zp7Hjz0EXQhhk7o7nNPuQ6/dgfyuB68LMr/wjtta2dnY/dOIbJzOHwsN5/iD
R+MXm+hXFiEGVk7Mq5ajs6YN2peBIbw3uVj0dmVNovd4mFzvXSsFK3QOJHzOwbFCuqZtKHEIUp9X
EWWbsjbSm9GLCkZ7inCD//W8bSnWSPFfb0P5ZbXXiUZNDrvdvBTDrrXR2miUhNIP4nPcYKyM3fPW
o7UOLIehNlPOcjHi4yOFBl40pfKgzEeayt3nDcP/p6sHvCNEtka16GzfpmI7QuBpMrdq86TQ1wBb
LDHm8TlQhgsOtgQXFjJaKCLI+y37dIm3pNqIvBRiemBJmYYjR4UIR/GH1Dufjfu81PRuRRtoSEtz
SoTeLC72b/JuBCHvoQdYIHpJMscF1V1eng2FplKfmeeS3mM+1khBSp4O4M2pgWmmX+aYMXU+1h1c
waW439U6peq3VCsHZUzNd3GBZzGBYlcFfT21nhY5IwCxdiHLkSVepchbVil2/jBg8iWXGc2rcrjs
QZj6AhVdjyqAuZQRYEQHEQ2ACTqGg2n7tuaHbBulj97p6pwMayPQlp5ejefLlq4v9WsXNzLoyPTf
x2qDPZYNamSC31DdmXoflQZ5/PeM7hd93W1sSDMWCUfeMgC4/tY1HJz8Ua7GCLSTjmSiS3KzgKch
FntER6VAGdh4oni+LGpqnG6YVrcfulYriKafGU5BJQZq0clVH2OjJW0sfDskxfICPco6AwEKcx2d
5dj7JKmVEMwfjK+tVyecoz89vFoNovRBPsxI3jektOo8NtZD7JYlsh+Ko8meOnjNrVPgcFvCo4yT
fnCwF7fsIJGHV+3S2IEXGxmDzVD0k5dqaOnr/S7jw1yGTwFmMVY7Pwerjv5q9XwlakB+LriPKvWP
y9vmeX0Gd1U+r07nF1hrJcgN9pMpJFyJ/ra/QEiSE+XvJc84uOsDIPaS7cZ3SMaaIBnaz5zf3zEU
z4NZLnsinzbXHilnZMNQeopXTag130a+mcczdAIfV+z8CFCb4QQARs8f2Ah8tsRo/Np/NwRpIcTP
p5MzFidrfZPY1BRO3LQB0Sh/IqItSXeEeqZO2vRXi0GpTQCOk5QCBV2q8kTuSvUXnBOU7Umv2Snh
d8qJ8NM9MLQdQTQkAO/MGgBP4LtaqCUmovcEaI/LLbVXpAdppAWgbYxCAmspbczOdQQ41sXBb8J5
Je5If88R+zhtylOCenTYCKy+ImbzVH5jUSgfgYTAVLdDLJ1OccwpL5OY0gPRE9Q6vNpeWkwcqjHq
xO1av+MVO9dvHbNbMtw6JGDnH4JuQH694NTYIy2NCwZWZOezLvaunCootQo5cIb5nK433QLfMLHK
URVoOUM+7zNOj/zYoIP+t1HYJUJy38gKvVpbNpMznXOdoQtmlkfCLzTWvqBofv2Iy4UmrzDjlPiZ
6Pajt5fqVQICpAP2DfHA3h8e5z8KmcryluuGBqAqtP6RMXxi4XYf+vaDaXySUJlQKvnyMAzS+3Y1
/wjEfMTuIqYlOXcdymbc1mmLI8zKxSATvd3juSzZ/3TT3rDw/rV5V/G0ZEQqSJLpyNRZBHT9Uf/3
mwepfPNH+FAmHHj1myAnPvMRBqS3duC/4QQ+G6rze3KNW60jbcSpiYNF11FVcQ9OiQmu9HXJ+Omv
oezjeRg3Hift8xjtNB2LH2ZnQcYyJDO6Iwz0C5A0zerd1DgNQu4w1q0iEtEUin8URcjRomH8FCMj
xX/JYSD5gqZ52Fk4I3UZy1OxBxvGzXL/oCRaki7OtSC60xMr9u4oXyyBPLlhJQm+FYFCM/UqrYjP
L3IOgQMlMQhG1LL1hTcQaY3+8SVrn7MylRwc7G+KvJi5Ci4C8lvJ0VnjkT9rcM/YBcGoDdQhz5U5
G9ovm+zm/7DxjaZXlv/9sJAGBqKgctnzETN5S+V9+LsJ7rLoDyWYCDXG6WWhgZuJqXFxLVKsEvD1
7F8DS4xcCXjMBU/hNBBu4wUpvpdWO6UTrjCnOQE5F/Ili7rj+58EjYYqtVQzaDOcaYmU2rRDlgM1
2PBbFXzx39RmeRCma0rAITq/CwG+7AVzEnuyc7cgAQD0whmJypTyZGziJVVk/pIgVSDGgTmrsi+v
9SzZ26Ctvvdsj8ugdgFVVugCDlZ4oNSXsamPRfkO9STchf9+0XAPlnyGElO0E5s77n3WiMxucyw4
CrI+B8jtgO/W4UiPTPMiYOLGFJQQMvkYKIOCaTclTv6gphmK55auIHwS+Zn1ajgVRWDOnEbTSZBw
9mElLKzawipCqD/2vBVxIa3oWFFmxjoT4jtSfFBGls5Dx0wy+xVObMCKgWvZtvJqpi9+urqiK/eL
7j3B3R+BSbzef9FtTxHxZLFYIxPdcMG+f+O743C+0eQzLwI5wsBu+qqh0irA/wjnkK/RPIDWSYRa
WZLRPsFiDdnD06teG937f1GugTU1DXaIP6XAi6RuSJR6uSolKWfhupYPiJ9bCEXhhZj/JaQ1ZZjf
PjzaO13XwBBPnCFwETnLE3b43iRqMI7BGZiv0N6dmZfKtREMEE3aOXUIxfXY+RRwM6DtsUQkbmN9
rpeSpOmFLwxYr3fQFpfh5aGllxCMkrxyhb2uT9QNxJ65jO5bxwT9AkkF2JfjLjBPyCKuP4MsBV+2
6wYOj/3H3VVUHM19iLhrHXQjgfKey4Hfn1IByIG6iW/f1msdby7UpzwBV8vanBqvM3JZuf+LBoRl
AaesN4TQJDbc4JA0uq4WzXcdMsapctgYnuz/kPGNFPnpVBQnX4UZTli16VdRL+lldaYCTt6dmwFM
1Yp/jP9jbsU/49YIAXZUESWKssn0lAiFIMsqtsInpjiDHhkqLzPOnTTna4olTYf1B9RfBQg3CcCM
ige+bfYkg/+HnzkzjU0V8BCS5sZtREaiftJvq5EsmRNTKf5dT4ggbbKySUM3aTfJk7U1byjXhHe3
SVGNbu6Xh/YQgSob9dsTrL0y3M8qyR833Ff4VIaN7VrCs7t2PgoHd3gLBF9Pb98xF9xQjXwBypKk
ZFecWFXnHmDx/N+6GWvhxumlxKwPohIMs9s0Cg8JzfOJ8U334goKofNMeJYWvj6gF8Hf5pS9senB
X0f5EGN43RyaTFjR/oG/SkhIdABhhFiqragerDD/vUPMy8rsVwMyI/hXkqT0TdHDnVRSa06xB+cL
kSvZ9zTW5jcSracDEfW5NCDOIRdyElB5VGa9I/kjDBFfuy6dED4CIi+A2uO6sD7bV8eJKLIJyTKN
QP4VW6spQppZGroJh+F4jD2d8xpPs1EjYh6j6mcAcLOGryg2d7UwO+d0gWEB+ahBZhNaCPCeUW5i
gyv45DCHqFPftdt5bxdGqjpAzbLhbBp34KViq5x+iH2bMawv+vCT00AwJG3oIpEJ/E7N9C/mX7kY
OHxdMvYLhVfKqnUge+CCDWCnRQq1BOvh1G62nL5m/lnyCLK31AtlpBh+rALHOcuWtfrtNX2+x6QZ
wzZ74vnvVlKepoTWdtOjHr7AqSRrIOle1uYUzeFP0ifidKgUTzXhSUaaxSOBZ6hiKiRP+GanRDoa
2P6LY0vQ+bQvfiE8bFeCruqfklEMrbTn/6Hw8PmbCktW+KNhbpa8pRhuL3y8nfXK9i521nwR84f1
VodeAU9evejP9bFP7JMiuX4k3hTiySNpzO/3S/ssQgB5AGXQohQvL6V8KJSSM+jUbBMp5T77Zlz9
Uml8mefo00dyfZFfsMEMrTy3GmMHHvpnQeC+udH+Md6QN76Q5lmUvl0RXgukgQCcvSYD988ZlaMK
rIZUW7hbt0LS4AvC/auJgZRhPcXDpb8zXiAc1cO9Y0pZvjh/8Ux+JmpwXGBUP7LXMgB/kxkbW2L2
sHgPXY19kZBvLSrx4WkBeuUdBYBpUZfPfG7i6i8f3DkLogyEQbwLJx9Q73uSGUQzF3iFNZ3AYvYJ
Ykr/mnGv8sHljCWPYAGu6JkwU+ZPMM2ypMyccJ4SWVT+1boB+XPBm1AqajUigJrPnXZ8qaB2jQhN
R1i5/OiUSzYxwPgRqWcgLHjUGrR7fs9QToLIe0+iSUM17BT4LKLAhAoj2RJLvQVO6ztEOmgkzQFj
IzqdhyJpOHo/YcbOHTlgh2wJi352kNfz5kcJUrn8foWWDgAyfjJtP9FhmQpf0wELabbref/hjFyv
TfMN8+qS1v7EKzVzEa0AD4rqHy9wdGjFygqJruwWPJLshHBur2DhghHBc/fWPYsNyrKo6IXnTZfQ
QtbxMDlutMSN75TNF0cyiqdaWgk5eLZvp11K6u6m8lp84kDkD/jd0O2MWEyUJkBEIFAf/S+kWnq9
SB+2bxvM3WNhmnFr94oKRFK/AAfsnWwCa+hw6dw4FBEvH2Vlr1vJm2QZFIW9d2Dw+EXxlrUy1zC6
SIJWOCYNglrWSn5s0unqV3blFO14yY8I57TPb0gdIa1pNy++8tK4kdTVliFm/Tmb37ITrh3br1V8
f8jQx4I9DBlx7AMZiyr2X+QnLc2yaKcJEWRYgNvWqhNS20eCjAqGZ2Tfr1caZy4YmkV8zhxMItou
pAFEBlKVzujNx/sAAq3HEdIJabOa/v/RiDTmJpijjhBLBS2bjhrjO8a21goc6MW4CMrB0zxjdNyH
YU8pf7fnsJdJ/y2KiixUa5ZIZ+JvUVTwmM0eFf4K9huJlYmNIgvxgx/Ou3X3kkFEu786tSQdNfGy
S/ALLR1dbefTwvoJykkpgnx/9GMY+bGBqFbWGOzZyXeDAEtdaptdVsZ7MwfzNJcsb3C16uSF1dTm
6MpYILl7vkNLNGCwNLfn8X4aX9iCk/ZtwaQ9WAkU/PL0/oiuE+urZl5wx/HaPIW0o6O9bh8yCc86
Qru8UeMCGkpio17eBsJjtHWpBX3yWWiRALB44grizP65g3BPQgfwI5syI1B7ZlfNtqGrY6MAeGTy
2ovDxEsgrfrFgOIHmR1dlf9UewDigoeNRWH6mpKB5gNmrJhzbn7DN3DEiAQWssMG2duV9//199NS
/vxW/XWQkkbv09AkHE90hq4S8zwLTqDfh1MwsCn9QVdgefPOALZywodDgKn0RMOEusp1O1eccQEQ
QkVynyLT0MGNImA0J4V3JTr3gNQwnmz8eiT9BZNrCnfIrklU8IbPAzWLEcmGQmuOZl4Y/G9SZtSx
+zgK53g+hgs5ff6cJyv6MYse53fCObTZjHxyxgAPQufq5lb1EF9dXH9rR2EnIzq1KXGn1NGbvO1V
vzz1Lpl9p1mHsQS8QsJ5uabnOZuQBlKTSHkJdec22B8tTO5II/rO8RvC+vCabyATtKucca5Le0Fr
PQIfDPGWLF11Gso3ZJcuXL/J4yfQQVfZekcmH7cJpvuba/0qubxR0ISAK3OgpCaJJpJNDE7Yt7PE
cDEYgSpwaACxpcmfbLnzEPsUYCTv7cvveUBSZEy2ZzwQMcBgKLuJv//O6kI+KNRY11gpfPbv8Rg1
iLbp2I9UIKkpbwJcJtTHKU3VbiycRuwrVXJ7Kj81x0LuMOYANLOgJLz96P3FE6U7Iq9UAbCW5NND
vQlcm1KMm+BKE99UG8nK97ttIOVngIECPV6/ls+qnZw0kxXBD56OVa+fd8Udl0pVjCfskFNSmd2L
T37KnnYp9qOz19vWK7SQnfiB+9kVkuwxEZuUbuclOhEevbQkCwmeHCSB3xMkHkhHEoR3GZQGnnpp
jZPuJTbv6ZANLzgruuBdK+KDNGbU9jHe3pSkfgSHo2HS10gzMLan/SVyRSWRr9HG1nTUyCzJlrxY
GbSmaphHYKC5xPJieqm/N5Aj3xjEfgDXVw93rZohBF6MRSugM7yH0TTIlKnxYRKQZeBbG2kz6D4R
kciQhnVxZK3xzXQDCjOGidmfdX7yVxXF5uNQ5K9lqrwgresptI9+8sTKxfEviymGlYfA7ANC2bfi
ajNXxC8XMLaGwxKEwihOEI4vl0wEft2kVMrH64pboWFJLjBEvjpBV6pV1gOzln8XOpQ+Qk61SEWk
GoHcr3zinW0PfskUQ1SnKlcb1hYrtIsIpxsIAepgY0DnyKBcJDLRzVlb0WLEUyflWrKok1XFAv6O
wWLLJO99RIreX6ax3L7Oz6PjTj2kDgc9xpU4br0fiNPUXNEq/xzwpWKcdnblSVr1PPAmYMy3Z3iQ
cA9RG3TJcWwy+5NcGv2l/BIQr0SqMpOD9PZMDlBSpuqMytyYxdan46/93boe0KMLIRAgacmIMKrT
7Ah5o2aBAhrSn/pSw/USyJAwp2O19XZv20yrnqxD6v2ddIOgtIrhkuO54uUY5x2gqDHLZ5/NRISK
mZCYpc8PpXsUaUSqefd3I+8WCvMngzXtjRmPGv1RKxZGWCSzx6FWpNJ9Tvi7RQGx1N8mCMaB297P
4we7vfdfLgbuflw1HFvD+wgZ7UuGeoc04yoC6C0VmiylOETeFWqqfKDH+LEgN14Dvd9ehLvn34zt
BDZtJxvznfDxXKO9JrFV8zOsUueWh5Fypvw40tuH1K0TqVWoK58d2mKdqOMwGAO31Gfpsm2Fc5kE
VNC62O0fj572GFMdoZ43yg+elVRRdfxogsD5NjPTPrjwqPquJnkNRGrF0FKJijXXwiBCb8oH9wQB
1JY+dzAfavJR0bRVYj72DmVYNdd1ISOAYDxyvbJYOaK4Nvkh3clzxlnj72RuP+ZE8ncSl9Ool4Hg
EvPuZyZUq5OL25hOtcmTlQ33aT+bDR/O0eh0WpyNbIowkqXA/dSFVxcHBwExj7VLdQMx0gsMe/A5
CduHGuURudu7B0mp3Ggj7Ck7/XHtbIZ+cGNCrRWgiH2A+lKrRs8ld0pLPFw2J+iOSJc9P3fqRXqg
+hLNRlHeaCeTzg/OK9/uvUBtnAlqmhQhucTLZs+auwyC7nHXyrhZu4/oxofqnwoxXMGJ2Dk5Bhb/
s0lde42qr2vid5edeiqahfGXBY6VBYu/Q22m7pnLzipyeL2onVBGzT1oPJuWVaQaKnQk0bWolOrM
kx7DqFU/L7csMyGODzJZNcdN6E+XyFr8J7U68OjF6RpfC+z5ZLonavdadzdD9BXUONK5MKLPKCll
5Qd+cJH8/2HBbBbZgAaJKZZuJi8HvKX48k05hK1vVrHveOPv6Q+CD+T0UGD1ykRJeQgEOO3RZVWT
639kwJorHnoHEGNTFgaXmeu2nmEhnbUDQgBkQz5cQYqCzbpH5RxCvqjK/otuhgbUk7XVNNHKIKa1
wg8cGyyXAcqlQEpk2wREdXKcCGD49Q0RoQdbYR0ITGFZaB8doPXkFqlG8PyKBTsnSsrNZlFVBOom
OC70wsNRFCON8XCdXoxoGxCEv5r9kipc1KDEBLD8VLLMw5PX/7KWBvQ44z2/mWjbpgHGbCIYnkkP
G5aeQiBX7vo2F62gdh4SN63EMj+PYKQmaRUAdLGHgVKataRhXDU5lV6dRggGVBstkCXwzBA1MhlK
pvPsnZqNiCI3S4Kbo6uBvkHdiZvkcjL6xzkfLzwpTffBSjdWlzJy8J5zkaxNVFLISMO0OTLq4gEG
gzYwWL8ovWoJFx7eDlmnpveVNu2JH/Tpn5RHK3TOOKWdeikAJ4amV3p5aqUsWsAYhSI+oPEAQk4I
tkBP/4yum5hUTldBF+3DxWTL6jvfpJ8064ufLMHJNe3K8H/tDWx0w9IbGV2O33Qa5SWT57aMjubP
10m+SWwDf4qxexSQzzlnQ7dTmILe7hXqyzM+AnrOs4et3Pb1Aw0Cp+fNInb26+UoNeBKFp5BWxUL
51MRtCGMQPXyAT7vxBWKdIad1psTruCCwzY77cN75PiqVYaDHgwczyizGgc2/7YLszjFvxSWDyLt
zDBsC/mMp9rVSaGr42wXqaJN3JDnHTGR9dLGfcjI6/ERkPrdJx+8JmBkLsfndyN/caSJVDthfLmR
yd5QG6KDao5CXt7FWK0gbNED9hhtVfMPM1PthbCE87D2bMbNodozzBsqgkKd6WdUfOCnhEWNTS4C
27lkz2JCVy01ZZk3Uyx+EVWh62lWaNIQ42JY+ROe2StDnCTrSw4/xNDcskKleTu812KSzOYHx8EE
xXkyi4BL+KEk6cquMn844QmqEHMAVgHr6wu4ZlrnOWrPPzq+6Y3ScJGY3FoFTxD50nF4zGfJAHLQ
m5EM4k9MTI+smcvy32VTfmYiZ53DQTFRCSxsebO8nPUPzinKESuYLS3ABI6NOkLER/Fc9lx+J12h
YO4iOB+5cdu3C1nkSdlaTi6rVC8m+/hp+Dy+xLSuJnUsRMImGrPxWbAa9fTs/wldul7s2N1XWJA8
3Fi0TVbM6TOLyWDRG9wUt7a+7KmT+OOvS+AN0eQ1ZJIqowE31FKrazVTVGJXLvlRkxSi+qLWt3bz
Ln3Z1U16zCn42CVJm9pM+ApTmQo/OZ63/LVR38YzlCyt9oycDIAJY6qevLAJqwsMmQRCmipQL14G
wgGuk7MPCKNqf1VuI4yosP4ONTdgbODQ8HeNi2daV8gfHT/eYRhMcfkbIa9oiVmfx0vKKppiAUkv
IRoEp6g0UIxf2zGMTqvz1T5XmeWzZ08DJRd71nfccQZ2CcM5ZR3e/ipmwiYRFLlWourPqavzBcIP
fw6fjNjipUhrB+pMwyEkZ36/tiXG/giOc8N7inEo1K3MMl52OQ+cOH0yiv5atyljFoo1RE8YbOrI
PJ0ZATPEAwcelrC4Ni/wobhpwBPeGW1PF8Ga1jwH/Pc5F34orkHSMktIqdOkPTv01d4J+FDPjl1u
q60QiLGRI5XyPCuSjo0I03PC45Z2udTzK6xbIQaBZbM37E6AqXQ0QNr6t/oCB5DY9sWJtdEgfIGu
X7L6eHy+h9EgtyM3JF7tIEOk5tE67J0H/vbsMKaMvYVslWeIVgV0lVLkSN/5m9kYAh8JRwayE9l2
XWkYnKgZb+R3YEba7QQ4YwekjHw+KjFTDTBoXU19nIvTyvBdKAx7l/4GEfVoJRLGR4uRVyzDiCnA
/1b/CwHNDEyKNhD50nUbPi5zMzvlDBLn83Pz0FTocHBbhOLQsWbN04wWCtcv/QGucbPNMHQkWWP8
c86UvVooN7jNp9IXL95GkhF69QilVHF3y7oo2/rdWOdCSbHvHdZiAS52nYKhovnfhibhvhG/Qd7F
zV8O6IpFfYPjn0IR//pILX4csvdgFy4/B5UAmvgNCe97D4L8U9+sPP5ZdDfS6wwr6pBQBrYEYx5w
kXDpr0TsGNUuO7QXtKjDaqfL7lPA/XkufhCt/JtoVJii1PpQ7HlOw4zJKP3MCY2ALljLyFj1W2OL
ZdSv3M2OjwyFk+6IrrlUUYFTjP8WlMfHuGGlR2xM7mMKVA4UxxeLxkgrs02v09tBTCvMGpXLZ1mR
et3EAuoCiWnbyPVjckSJHgGarjUCn0LVCbeex4bSewQDkgTcf9Tb1CduLFhGUHFUJWmIeBdnVHGX
R4oobn2evUDFnLoaFHD8UQUm9PdiqWheZEqUoHm2gHPobkiPJtpKDLC5cEaonlRccxRb9om7mKNJ
1FmR0Yqs7slmXIOdcQ2U3amNsecm3020QacaG0NXWPig8Q0QuPW3hI3nBEqw5yH2G0Iluygyxg9U
hVVaINFFk5iAkPqkv6ys1Z624S59yZ8T07//nX+dVOUwPM3gOCBetzv/OE2uwegfWk9RmtQJcXyD
UNBDksm/yAqcYTh+EsaK3EsHvpEQSkxHfIsNSvetEN2weTH4vW9BthgrCzhTLPHfSaGVeT12E1Gf
38e5pyfiyWQ7JfE17s8qIj8Gkdt7vA3lnXqgdHG5iqws5xx6eI4lZ1kTzl4wxxW3BdLarttoKpcy
97jIQa7hRVyMrREh5Ox4XiiUZ/Uk6UZdtLu8503yJhrcKRr3AXhmDZ+dfV8BN01pV55fIXW+UN6C
hgYVNs1/euLMV/3wdjJliMk1/OO3xRLe5k8OCU+CkfWib4E4EQoIU64M+g3KVd7od/ooJgPWZBl/
JbW1MoqDeKfPerUbI3extDZol/0nZmE2GCYzFoM0qIVO7ik3i1NPitLhoYnPl9guKBb8BDxd5bp+
26yZAtWJDkKXLKcphBMtobWnW2qGuMtWCKmH3LXPPVryiSeUylJ3xrvL2cxCj+iDJ/ZazrrWCwxq
iHQHdX0ldYwVI8AcPp8UY7wY98TkIoMTn0DH2EvWcJDOdWIZp5/u5fHXLPHTexZymJN4YQh2aiQg
ZhQ91i6puLmNS/HeZNAJCZyo+3aB4d9UG1j5PcRzPUlHI8GfXsaSVTydST/ViAyE0k77H+wkcx8g
ZQwOSCxHGsmOXuuRKITlepY+2qGD3N1veaINmTf88a4yqxo5losXBTKOL9L6ew1ewQuHWSJh5gp2
tnaBCrU8Mi1NcrB8ODXpOJcltTJRluBO3r4fCIMCLgYsA2C9a2KnGzv8WbbSyLIJmQQlR3uidIoX
85DrGPaidtJtU9tjmEtuZE8bkcpe54xZsSaJ4iiLIwz7nE8dKfDNf08jFaNi94VJrh9duLXX4Yel
UC805Q8nxRY0qkfwNwY4l2f1KY/L38RgJrco8B5sqkD0aNQY1wu7Bk2RIdj6uDrxm92e9siSqkZf
9alF/xOOp1TRDjQl8tHJTyoW3DlCFgzNi5ojVL4AVBMGdpk3Ue7ZgNuywOHQOnzpk2t8PTA08b6X
dE903RHVXmxC1E+oX2Dly1wpkMGrkNev7ZPBwaXcdsRk2q+8O1tXY2zDvvo3D7o94L175rQXamkU
W1b9mdcZkVfYvSIoKTBX2iwtyZZGrgpfL+jH8HBdz2AxRk1txZqKijs14m5Xds4Y0ocNWAyJRGEn
2+4Mm3HDm20CaEXvfuiGpkx+XwzNEiA70j3drzCFpxT+do6Q7XrG+bRNK1rJNFYDbbHIhhEcS0UH
dYpGLuycZl1QU5DEbfzYKKSQzFsMlS40fsC0cUMnP4j3zhys8BAWeyDuA0UemtIs0KgDSmU7Hxck
cUxv/2e3njlla3ZgksO+YgGGDEUpU2tsKbzsudIIekwoKzfq9jyoaOAKX1oRzOPhWlEFfWTpj5FR
ytLR6r7yzjFSD+ImmMX5eST+LX+oPSv+pvQgI0PClxqg+Ws3/Do4NJRUcLo1zREOSQPIN2fc6OLG
156cdisNdpBS8agi+UB29CgzZP49wggFrzI36F6M8jHz3aJ/KvPbf+Nssv/dlupeAoQe2gMQw57w
Mwx1IzBb6QiQNq9LNnDGTbhy8UfqqegSJsEh32/u99AQYaAz8ChZ4RnRF6B1N8O7Xb2eX+bAXrw1
1jmTOMcJYGhApYlUJfL3nQcJ9bdnOBYJXOrxuSGnsjDThTrvib6z8L9QKN7td8yzVCxUJQHKZuwX
SNVCb8OkagUJeGVCbtJqve2aZQnFS/0km3dH0IoLMfnz3RtpYbGdj49ndutMDLMPbSdW5R/9rM9o
rflnDZ9Rycn5Orb1SS1IimZW+vvlrBF4QZlFjKar6odhUQ3+WOIr7qajS0c27KwJwIvYU5ReWCWd
wqL2fAI9Yl1KmSQbbXzaznopgmB3+p+VweuaO54jTs+xCy1Qx5jWB0sOUsY5MULk1f6KTyfdXAV3
eFcJ/urKNb+lwW04WC5wd08wFC77pBbcFfR11+aToC3kkjzPgCSWMzfjfAgMqLKR+E2hTLC1169h
MnF+Y4GIfPP9kCe6GlP9jUj5A8irKtAWlyGk6FPeUQI8EGkHqGTmb5ShcSZGSSLdDZi9gCByPeKb
ucJ23UUqnijb98yZSOaoK3qYh53ijSYRHCIrC+6mafgAPBRV1nPEOBHA308BH0M/LrI/l/L5p+k7
ZeudUwAPPlhic/va4i2kMhAQZS+0pUkmgLKx6VU1q3UOZhxsWLghExFuFrEkSUD5fFVl3AYk41Z7
o9knN74E3lUsijf+ztoJ1hP/ndx7HrM6VDOdxjlQjLP7BJxxJUUJCFKaZV5VHgrCr5uxKNKgeDfh
jS5BPvOgHjh8XFHLlikNzZJfLNlOFKqo0OUZA3XmAmhfw4nYpuqzBuDVjmLi4KyASGx7eUNqd5IY
LNSwrYbSunVBuK9KkPMFgAwYlZhw5BQla2pDic4SyfhlztjOoggPwfMmR7tv+7BJ2CPldCG3veeI
K9fl34uQXZ7/uCkc5LbvaVoQuYp97jW7CnfFKsEWvJAzYziD/K7E8WnlHI7j6Bu5rJWJLdsrsPmu
YJQIMzqGQqcvwKJsjIl5Ouz5VUjKssFYU4clpaKcMTjEEAmGLooluaj7LhSBOtykYmH6OwNeKtlC
MI3aAWW/SwWCENxYV0z0nwXB/CQlIryszpONCTLTAj8zNSOIVomSwmu8ErnEHmi6ML9rXSrKBYOB
Sj5qzpK1gV/z+phwS1kSIVsDTRP5jz1DWKK73BpRMJlDFWrvWKlrBbvlDkYAPOYnRpd+lJLG1IXu
EfMh/yEbvTRUBwzPVvxdc1Vj7mJpclcNgleUwCidicjPNK04GvV0Uud+Cea7biRS7iPON6zLPUo+
WA3cVMDYDB8seP/qnAXN+4fhzN+HkUeCGfLe363z+yQPmolToB5GMNPCSv0qcPyKysba9CWhG7dj
20tOHOGpRlEyM+Iy6fGt4/MiZwXAnsP3CAf3+jiv2bShHLG8jKRhajH8Vn9XPbuSn7DvqN7D192g
RJBxwNGUVqjFnD6Sydrov+yPGLLvJASZoEqgUhGQ72KZSAQDV3SAMAnaWu5KQg8TA8OcLEgwxgia
+K4sR7uz77sUIdvwcDcaxBdenDSJypIdiZbA+egJXQhapTGSmQcfyu6vbo8MszRi6tHDqXVN7uM8
//M0S9xGxZbXjA6jD1v5ypeKSSY/aDt7aMZ3vBjphjhScLsaqLNmw2mbssemzstUfHwp0WjCtygl
3UfkiiZlpPUoURSoedm/Fci25l7EE60Z8451XVIM1BucMAm/sFMO6DZsjnQa/hpyD5Z2G6UO6p6L
2bbFRN6UeffHFK9tOcSOHwwV6O1pmuSLsrqI5lniqWFK44KTLwK+CCSh6mHiN3tiHzryAvb28K3h
G0u1b5R0mke22W9uHwhGu2DBFuknTowFOAQ6FdWdNr8LXTv0CwTheAYG3csJfkGT0wiGip+XDCtE
Jb/E8BepS74hpMdR8kov12x9VijS2WCMoCo7rSs8S/RWYJZRXMxZbzKpjKrO6IeT9XwPLOBdlaEQ
VcwPHcWYRYohSkSArFGj15GEdLzWS5nCaikJ8tZCPcvg8Li6iZ5pT7mOQQqKpJUXx1I4Iy+Pde1U
jhEkc2RF/RultYhmSiDI5ZVHrxEb85bitbRY2DyFNJuZpzWP8CuHo42zMExpo0qJR2QmxXyULkTi
RaoqVCEPTNk8JOzYaHTM0llzZGhc58VGVCr9tyR2GeWjX1DUG22dZW49M3ugFt5w8n7jZ5NqlGKa
KYnsB0WwC3WpOMZPsgvd1DoEcE3IZkLbXrx6CjFUXlp2bJnMmn9B7Cm7ym1rBMnqGgVxDJtSZrxn
J90mO5nvnnDUcGghbplGap2e0ZVIjtmfxhi9vyDIAF8gqx/7l2E/4eow+f8cbQZuEgjCgLfkNuo5
uxLQmL3xMFW1L3jZBQ+kbgIlOZzMSgR5Gd9+tl6YS6WPaNysNLnr5hR/HkYsbU/kmWL/sb0VGB/C
FjIPd/PclxX3c1Wsu16RGib6iQVnDthcbyCcKdeh9NLG1moC1RDKaair1eUK7AIbUOy+9V8HaQU/
/px2LFFq7PvJYpTMBSfC73fdfffDGHk6l4i5KQc6DlgxPQiL1sgzkp+TrtxjNeIIA+WfvwV0d18m
+1Ccax64iARCO0wwh6xTznRSlIczjarXRxkVGIOVZX22s0GrVGFeESo8908pFUaz9zKTGqIzL9qs
ibZG3vdffzrxZ6neV/dhzFRgnktstTqKc/xzzKonQJSxGDB/ZlEg9ld2SCv3cse41t+YZ1GnqrWo
1l9sgfTNNxJD5TgZItNLQ6+AqwXZ8VeupR6/17dGqOX6AwIiDLmWGlHs+IQb3qImq9PmUZaZoyu2
1b0Sf3sSrC3bgL7ymceElD+lH0XqGG4DyAnEgRjSrjxwHnOQ4nor5kDFWOR9qy9Wd9DmT/EcoiNP
9dACS0GXIx5MsptsaKA+6i3l9yHWwtv6H9QRnea32D+mohDjPoqeDotqyn853fOU3gVV3eiAYEEW
kqfALQKebn0J2InL/j5WigLXiomoBf+Uku/LVhrpkbGbQvVsLgGMwws23idnbPpvDi/AjTmRo0zs
0qNpgdpYdF+cmsrDps8pm7GA4LxsgeQoliKflCMhQhJIN+L/WYcunUUw0JfgmCe0xTk2c20XI/Nj
a1XyZdeCo2zgGVg0HZsfhJ1cJ9IqcwBqnzFW3L0dINgt1fXoNcxLN8At8k1abW7pRIKJPv4fVQ03
dt1/pKUiDST7+BSuB17eyj8LoEg8YUE4VvkZfHMBYuDs3lUM020LmQC7LobHk7VkYoTY3hjL1SK0
/ykqfarACg7/JpLv93LY9I4IobQmsgtkFueYiiAYlN2EKeyAMyba7n3bb2h5d1GtOEmucrUYBRjf
HY7Gk2Ls5qM42NRk4QM+FzkrzhaSuurPIIQQ3pypQmEy4S3coT2WxhVs3KMMxl7RGxK6gIWnYWMU
GliIWjXTM21wNXDzbfO1vlCoRSUaO0IEfnIVnt9tlqnJEvMYNAAucvSAXe1h/3LHVl2EP7/iDuTO
kCrLRLNFGquEVTTcJSoRrpahge3ZLeEmk0ZBJZvzp5NKjrPXFMYhb6wVvRfx/JLnK267AgMNfxzh
peXxGfOuF5LyIsLc4WkUomiW9aR++jzx82NrqtEc1HljPdpaKqyLgYkTX9jy3IyzbRCCLSD31+g4
Gt+jLqOsSQPvA5CdQZ3rruOTJibAfYpBekfkeNUZhkb18gHSXCZCCwWjKv7hUyqDoTWJFf5in/Uk
DeYlMqUedOe2y8hGIB0oQvJUjNdbkepFBMuWTOMItOvl0uC3RY+/cm861oUCC84I//KnFnxnohyQ
alokDotXDUBmoay1fpRNbE15z7IU62NNLKfoXKTdwuGV50FblpTh5otuBKmzysD6WlAy0KGnCuJM
tSwIurTz5cVRDmmHV+BCjAW2QfVcELeE/Kf3KWpoezlFePu8zJpQ/n3ripc7AXrAT59ZFKo02r0U
qMvvQwf09TTEDhN9v8BDh6pv9agtxa0RqI8onjv8e4+9m2neGh62+UhV1Jj44G+hBY+pRkaRGhSa
RjPL+f1e/0+TBai6uvpoCCY4R0LHhLNVNrxKJSy6pfRsa9CEVKpm1VyT3eKrOF0jYdzp2EM5aWJ2
Vv4KAMRlWmFX6CyFJcTyTri09xgMnOk1PM82usg5zyR8lwnORTvHEztLTb2J7GEeyPfkuzEkqfrs
8DY9ZJ9kulaijfjMvRmIwugak4pGNCZScYUNULuUIBgKtQNUOBPEjDGfLB/ueALZ/TsjgjumMP8m
xforallAX6fcJ5DNmhj4Ha+6C7pNqSJjn57nGIgr0cn8GjiWNXcEhZML6X6/FUhmQTO6qa8srmpk
uge2EivB1TzGXdK4utsU6yhOCotxTcUQtwnc+XLX2gdkhTmFZ3cey8H8kPsDNCjC23Af+6QqdW6Y
hmX7GYC4Vg5DTvlQIyN1KQF57MdXlT+ZNda8VIH9wBASSp6Dvvkcc8P1QrgybwKJpyzOf6Fp+Rub
ZDnA/frNjXAmYjw9Rj0ruK03ddlpcaHX50rA+iLyOAZOTBBjtEoaJ6Ts18cSG/bWca3NYn/Zl6d4
H+GOa8km2T7h5UB13YLCBrcf67JwuNLv2ky5skh6ngvaY/Zwbe4lTOvkigjEXVaphqn5pmKgxQbM
hwPdTgjJ4R9Behtz2ZBMxtgsSDo2nBFKpjq60OenmpCfrfDb+LY7Pqx2/Rm6jmzswgyIPw5M+dtq
cH4WLiv8OWRX7aGuResvkwiKf0Xd9sJ3BKY/bndFo/iuPsv/HrP42UK764THlNiQUT4PwqP/oOIK
NHJSHhRGDqEjmd2Z2Ku8lOaSJwN2ucclaaLGV6sehgzCW69YXdh0y6aV6YzJFNbgVvatyfo71Mlw
duHD2rAf+2/zangdh/50IafNTkFQPjichOaoqk8LLYsj+7DwpQ64qvBzZ4B79z742Y6LwCAdL+rP
IK8KTu43xO/lrfZBZkgEXdj9VLU7ckqyR6o/4apB8UytGdfknx0nxE5VLgGAyoUOMkdi/+npXzlF
uqyOiG7jTjtfKSXwklGnb+dG85i8ntctXQwRmHbQo6CxQcUlpGQp/YNcmODliY/Fx1vYGQzTALHQ
rl86YyiNgQsqxFPcE3mxeywHTFUQOSLRSlfJ78HA1jYJKE/lRmc9rj62ZzZjmLNTZpuGt/UhbRij
SYk6XOBjEBazbpDmz12y0UsmQno71s+3xg/uCkatEmtvEFaMFayP3L86lbwr+/oNW78weKZxTHgX
DsgNrkAg6rpFuwf0H3sbA/oyakT8eKQQMFBpATavhiOLjFt/zCQnzrZngosCDZnpjCERc3+NB2hu
fzzwtDEsVVFHZK8tp/Td/CtnbQBKbwrIn6IWv2tvGWERqqlgV4L6yDyccgWD3X0Lm0v98dn6ny+n
J58/FG4oyzbmqV2ZXOkweHCZdj7VNIQI0yGfoWSs5OoP3bTMHZycZo3XMBES4LSe4xIYKd7FX0HB
JZXDKFCtRfYjstaC6IfW3pWOSWtTokTSIeC1wkXlUxxBhe9ehu5FrucSb/gsos0BfB30eRmi/GMj
N2ctM1Y6rfLborsJlSE9gTygS9Cdo4ZkssSO0x+rPa1v1zadG2aJqnv4wx+AtcvUvti5Q4PgXHZZ
xdUDSsZZSKdmcURFOQSl24V8Ig4waDG63of6eGqIjiCX9GhjCcCd3Xxz5sOjVR8PdQcf4CA32asL
3BgzFCPLN8SAH0eGb3cHiBD6bN6fIDltJQadzcSzWZ3cqrFGO+9cVFWLfDaJzUIIt3DNQwLPyfXK
l/MIfNtWfyugxMgZwM1zpyL+oQJqgNy4eoaS/8PLlM+fY4CNAYgVS1F51l+cdihe5s1ERoI4LaeF
RYFnm1ouljEHjcuOCL0ZsxeMfuKvgM7uOLEI0R669+3TkPVbmR8rqH3/hHrUYzXs9OIp+VydDw7j
r16vH0jfmX7R2+3LdbB0G/Gj3febkQRmkU28d0kzmcL3u5k+mNCuMTGz6GEKj9ScncrdtUmq7C1Z
R82fRqW2ifQxKnjZ0uGuO2/CF/w9yxnoFMpgLBWr7xrfRtHq54kzHsjgHE8ADjriaUjdXEX0omF3
uiqwqDVDVauBj+1/rwhKh0gGBhs2yhvAWg4cdAXp1u6ZsSEie3p7a1KgAIApiXT5nYOiK0SvbV9P
oihZN/X5Uklf6U/3IkOGdscGeG2PdpeFig2mlNbQQpvxYQsdab42NYXfWGf8F+i/Jh5W+SyfjgUD
OXzHYZuvSLJVLoMW4cYgxTF8vnFhvecULaoxoIC8F6D0WWM4fbWncr5qMKM10oXXahdm2jrzKaSH
RNanJ990nGYEF+rgjR+9E740t9m/2mFSRKhqeeeS4lC9VOkD23jJDG880B1a/0vMN8+9ubAAoMfJ
cHquq1SQqV0WC5xD+dePRSxxVAuuW+7weCczS0sedaTgMv65Z8CJ6Ul27Ll47DklOwO0K1LGhVye
phkxB9rKxfy1KI2F5otkIuGI04IGoiEwMZ2ExoYKzYkUhNo+9pExFzXcni0VVhjlxCUIOG7NPZmL
D1dElWAwdsGKtjnM1/1GgevEjjqURRkO1qy0DEZ3dUlixWt5RreO+OJMjJJm6Dz32heed70+5lYb
GAFRnVWwl14yCGQ1V25zsEEXL9UlnrmK4wiKg7Xje7/jaupUejBDCnpP2HB+Di4IoUuQq1SlVOM9
g226esOTf4LWAgGCEjad4AlBrfd6l+scoKLc21298qcEHJ9Rv8AyV6rw9Ahq7KD58/ozSPGfmKnl
xHkOGkBGqY0GlCVLHL36z/blkDTDOE9ZdhlXLNH8xvobhXCZPUjOVkTEbuFXYQBP70rjQLJEi0CP
c6slcPu8Dm/HPvLMmNjpOoT6Nm5crxo6WcV+Wxj8sOb24lDKGmvKVGk1vE+KRTLE6IzSLGRAuObE
Gx0vtLOXkIQWNQzPe+Vx/51bBbNDtCe7xp/kQ1J8FuyK/Fg6yp2Kym5FpOwGbksm15yvFpckJhOD
hhk3JceyG6aUGC22AhqLB+aht8eSEbw/qjwbHz/zIRdVXWnULVPM90Or7mdCJvzpd3IPqgLOTjOs
ZRpnETA23Y4xGEYxPOOIk/KHygHfNh5J6NwrnUNDdUy6oKskX1MO3veh9Lb6XA7u80mPEWYpwSpi
Pl1/2gwadf/mDK2xXRyWvChj0V0onuIr1+j84Bt2SI3qX8igTvms818diXo8eZA4Y+IcZI//NnQc
Af1ENdu/VMwVrO7vU2MlBlPvD/ATuhgwaJPJTqkb40UMWXveSBlPpWeyg7it86+3FlRtVfOi47CT
YoWSoXgKRBloycEwc4K/MIdw/DewgS5l/WbBKMcms4C2Kvk1AsOEFCb78tbKxfCOX1Uk1u10WCB/
HpWDp8MS2JZMGb0tSyJZQpplmfkb7Itq8kX6n85dRTiZj3nvqznxOLf5U2gvbnkLsOuPwWLBnBrf
FNg4cdAuHQJ53A6wC8qK8Ju7wfi9eVeiRcFYozh+9h22KE2YxplsgfjMJyEsYQdsq5f07vp0985B
4zqlU5Lm48dXRu+OvJDocvSPjUdxrSgdeCaIGwrqFnzdhtXg7ostvgAK89At0gjgy36DdApovbMY
bTOgIwid0CPAkTuBlZYKJEvAHKbpmTMvbHiyWlC+iAY+ZlMIU72wDiTyNiltzXLLA7Bw/h0GhVU8
Dg/A3R5Ica/kdqCIpKjoOdvR3VgM4I9YBp277qTNTPe2vwzKwWgHydvekGgN4SQOMXNFgDeR9PIa
fx9K0TZRNMYt0kS17Fafa+72MMUwfNmW8bLCWNKt62bPcuDQWAtr8JyFyv+q4pZugdTGZZSu09Ru
4Q1TTnflgqXG+Vl35+vHhQFisC9iuzkSLPw4dClIwYTqcXa06SEugDcsbLtkc/wPsF3iN8Khpx9X
Vr8p0SHh7A5vuZYbYmWzwMqDgqshDgzCWxyKkykoRVos5I806rkqvo6fMHhs6mnQ1jb8D0SKCQ+v
3FOucPaWEyASMk3w6WsioweikmyTAp9EwhGcSJasKdzyP2yzfPhMULWUmWCMf8g3BMjhlHlNp0M2
LIW7ayl2X05P2az04LhhRIGmg89shWIDqQ+iVFhfC+9TzHIgl+L/iCZzOBzq6TvlNsYSEvwZBAGd
+9HnV9NsK0dIAo0/j4xk9mv5LU1zAMpiAzjCcxL0QdXBJnB/+bWufogSPXZ+EtmDfbvQp74m25zO
6+327ODQK6WeFHXKRb6RfNrIMf9u91nHYPzu4uHfdTIQvhDAM1FLG+ikKxHU+OYXAuxZSs1PZyzV
AFf1oEfnGQyqeTXlayQeUHm72JI9Q/RjfbZazD7ykAWirnK7OAEv1jJzZdRqZ0YF+9rQi/FAkzvf
N6EuAbPZJaNVwfoLJLuhepra9Ypm42jrk75m0b1YrxGTtImygqRuwVi1crEATaz4PleB/rKFkTsE
VMimb8rzG9fi9bdpujcqlmj+MOMv1F/34gm+f592P3NxUyIG+KMzVSk60k29jE6lxliEIkK0Bn6S
Z9XVLZLh3svSyMmYtv95gH6PCAbh3M3NLu6LHBHlHs4EV6LfBsEKJg0EazbZELBY7kGzwXY2ndBS
KhX0K2vVX8Gk24H3Np11pRG71O7zEYO6K/iYXd8GFYlL/pqtfjy/hrC6h0/ox26NrSWwPPFgrOsS
MhcefE30twROOwbTiwJ28bPRCaofaSNUjVweHaPPoHv1PSU4/5HRs2K/nhhSP9lQZ3j1Y6OIMfxa
xOAuHqTWJQKKrnB6V+ULK6vm2reQ5z7aLc4mck6KgB+orfJYUM8DrbzYXXs4E/ThJeyWrwLKvOES
2xXW15L8hZWaxk+c/ue8XMTZDjrxDe6x5KPIKZMr7hU5o8iw+NP9GsDae0jwNdE0xntNph/vQULb
1YHpixKO7+nUbov7lcDRnwBG44NDvqKfCcWJSzoLEeoiJAPr7fJMhbMTji2AZ9METxPRpq0sX8tg
/buwvyBZ2v1dCGr0IiZBG2ivNK6OblYYWvXJWFxFSzX1OSktgsxpGl1D0tQmfYF2iPSjxKIVJSAe
c0DvM2HIzjpuhSsCUsCtY+wNpjtXpIX1ryaZY/cv2BZQXFjrNjXPQLZMxOE18zs+d6syho8EjhL6
jYDsBDsseoe53X+Q4fvDPre38xYpOGJGnOf/2Xa9UXEiJEGCCl7jOUwv4YwD8k4Z32OKz2xpNO0w
8JyA88lrEVIYPLKAUvKePGF5Ts6d6MO5Pdu9OZZXrq7HFL9kPdrNobGYhTc+JpYPPRD971niVSpR
1SQDTc/S7C3fl9G45EZkSjC4q4yaScyzdwHf1Zg3uxm58BfAAJolGj3ZG2JhUdvytKwcJKmPk8cB
qkwmLcbIGpoEhMESwMn4QsaFE00uoOpupfKYMDK2KOBUB5NTgJAMsyaCTpR8yH2S1h34oz7Tet6W
9MaMbNdU/vbpneC3n1+cxKhcaBb/s0l7A/m/2QDgzInAUHVCntkZ/xVz37UAqtkqNtBUtxDfn/L0
tbXAmkQEytJz5y78NYIWXMy6EF7aWRG97p8tMCj/cnYjArC47fpjD4Bj0sL6CyFsZ4e4a4DU6YCD
JK54ErCRj7btBvRd23O/ZLEqGe/AZyAxXUhhjlODF/zo7g+3dVA+BCT03WNnnanKH2qjIziAbZDP
TOri+8kmt4thltw9i2hNA32oZfxryECC+yktnbveJ2SBDBFIdYHItFYBe6BktvpI1xlC/yfWMes3
aQpk5DVP4+xgW9b87WwXnx3oCPe5XtNqy5jK8y6NJtt3Vpiy5axfIkEzvYncO3yiN+x5SQ9qvyKq
y2Z5XvLYYoT22bMLMT5gNsJr03MyM9sWXLfyrnG44YyzJXu31wV0iNCy3UTTeciwNSwiKINrMb0t
So8R/05oDK1yisj4SL0R4PtBR1qOIkp/na/3HA1CbqQqQvzVZzrUGX6e69eTAKB1THSUy77JG5qW
DNCTCAiGtcow+KwXDRKVP0GHxLAHmB37LYZYQgK4K/IDCN+5knnieJxJufGU9UhtXCkym3M0mCQV
0GURIYkQ0JyF320VDgKCj3f2rjZTbywX08J7/mXPthF9PXDw1qtzroORU5qTAfoGrc1BIvbL3Rxf
BdQv++8paxh3d27jz9KYkK/FpXE+6DD4h6V2PNd2hH9ScKOdLX+xiv3toNqv1RPnd8iT6UodsFVU
IVg/mmSwg9f402kkSmtxSNdWHLrFloljsGiGnWGohCxy5uNlKJ4emPPSanS5JI1IcEh2Gj8oUmoY
pL7ZaOFy1lVwoSayYpwYuy0Hds8d1W7NYfj+Yt+PlKzHmOsIw3PLsSIFyLoWjk3NyT+KqDpXPRdM
nv2/3hQYNQBE0S7/j/A3TDV5D+kCeadtCnz8Zwt+7wUOh/M1omSEt/aaJ2Vcv1R6+xtBdbTWhMiT
2ZhOgbf9k8yek5o+9h54MAsB0LeQpsz+8td/+thiCJjw1H0LLWB7f79AVQkAq3b/Avi2brx+AdY5
Uomkzg+gwd13AbjjQ8EYrYV6P8XBjUHCdrtY/xKez+QxyU6DS3/JxFxuwG+FXxv9fkTZQZBSVnpH
oB3H3X7iH8dNpIUmwncIrMpZ7zJwIJpwJh6JOXw1OIu7E2nfQvufQ1RUw4KbIaoMI+zF3w+0akks
oUhzrDWrF6QrDZSgWisH3E1+nb9zB38X9GBhQCzsJL8bheZmnFV4MM40jMcpeNJxwtC+w/s7qAdL
bny372C+cgXcEvWJxYe0NQCYcac0s9No5qKiu52K5tEjNUCi9euE6rh2VHekKRAViNfGwt2BvETl
ZbxTT+c9VRzacVsMTGZRqZKHI0w7TKfmNs6WxAGL/QLv7W0BIrBrTR+TtYPwbNh0/hPDH6i8na7c
iIOQ4ADEGWJKqYeh2ZsirBwCAjOjtQvVy3VF0iNFcJrnwif8ViRtrx9Ru8iuKCZBBbH8vIJ7ON9s
sPv7s796gUOLFntMzvUG3gYxKaJdakMGlMRawB56rD9x1XH04zvlnv1GPZnYtRz215faqfNXdiYr
hEO/4B24pvSu9OsPfe+NbC5iLJ3MvKwG/WAsWIn2viA4tv0LWR3zRl+3au6yLtCth02zz15K2XyG
qNIH6va+xgSwoOr4JHsSTV/CaAwD+Nul5UoXzOxE+DAR5pk4F/2/qOfK1V08kU92e2F0iOyvT5kt
tnK6MbX9gkZH6QCsUtPYXzfNFanb1+IN2iUA0Q4EyJGVomOPs0mKPOm+PJCTiR+lc2xmmvKhU0Lo
JXw8y7B1iCoPzmAuZNuhhDqxTchu+6J7v91tipZ+G5B7ItJz7NTVewXypkXY64jwN0rDRGW+UvA0
UcvfpEe8qTkLkOUVPx37wC2oyVWvCzBAJdHsfgSTgpvCSjnWEpeUw05qRPxarwzgBgTFXM+C16nW
Pt9HHSEuPx1V4y/Y2EkgbNFzpEU1MOCMBV7go2QqnStM7oDYVfmqF3TwjX3cX+2OgdF5KHIgajuG
YEYrRDNFsxl5jZQhZMXHnQ7Vcl4y3eN5t2o+2nYszIl1FDG2X8YsTYqV7L5BAVpt12+X0OLkuXwp
dwomh9KgJZmiHvcllwqxPjadfpnydkWoq6i25wkgX2Ie126xI9tMA4NiXnxPTmSvSE6PhP1jPNHa
Hb+unDkzvF9+eE7CCjbuEhqotgWLIQa8+jLTm3Qtcww5pz6Paj8xLP35GLqZiR3lIdihjtyWyOvF
Q8s6A36YyCKftXzA6RRdhP0vQwCwpiNK7dICegxHhkiYNWonmdlV1e5tUNPu5CZ+3AsCgRu9qI0r
w6dF97rFY25b8nucbKFSGNVTdhxA91o1hDtSoiDF4FehhOb4gDulPP0F2d95FO98ycpk3S2DGpXK
ShN74/wXuYg8+V8q6HHc8hHl/fDxJGYNcDoGyubboNdTyomk94qGw7GzN8h93G4w9bVBEro1FP6B
WNBKgAwHUZUS2KQSoHCbQ7HnErYu5M1GLAMNqaGIi1seBdJ0Tgorrk3j7051p6o5MPLQfJmqxdaD
rsNw0Z8HkJUEtgRWLhBUNSK7oEz0CvMWIii7CudGNnX/JQETSn4fSxO5A9Breq+vjwxb4DWKgj+V
BOFFgn4aDcIvpsqdqnFjVqXU+4m3L3f0OYv/0Yi8Iy+ZQUTl4vq/6KsQw/p91T4CP9C5ET9UgmCC
j/cIOT/Jd+nmyA27JVEHSbgEfSeYm1WP/43DYN62FpTpoxtG7poCldiFP07KuLdbm9a7OnHF9AAI
OmcDOd1r5a6YrpFIeSPV5Lo4JTyakUONLMq7zstMz3kxAhtJ2SxCZWVZP+tkpcA3GeCwTntdQ1qE
0rijVRF2yVbf+XM8f4aGJdRZSPzaTJBOYG8++1USsZV0phiGI2SupipnFR+g0+q9oHsQGTZGanpk
bctoniQQAL3A7mpNt5L/gbEfMb5lf7pbZp2qZToeyo23etxixSbFMqehDFgDdVxfBy3UVhY6shJz
Cr15fNJP/x+QqbbtuVocb0eAMBvyEqw5vIGSQVkhaYcguSPRRIVT542/4ENIIH7KtjQ0YWKr18KP
YK9K//FJDDFpH7wbZ9moqJ0xtnZc1Rq5eVkLU3Wtc30e3Tx/5M8hoMbX8+pUytyrxwyMKbR2Nmyo
megY9H00ikUWPVznOqKMN1dqwfbCsWpYE7bbk/+nkabiHqtL9DvXvI7kBwTyJQpotv9/ozTL/R3/
D+msMe6y7DGX3Kzh68G3yjQM5N8o4e/bkbJDfWO2AXYbLIGvtOvGk+3qvUAdiDOEs4j1Ui6hCSwp
Pgy5MmsMXvHmwQq0XgkFw9N9F1C1KIxTXON7bkygzOS0u/muH5a5bVvjcBgy9ShKo/mRo8rvbpXQ
R/RytA/PwLVkKqszr4xvXr+Sm54zNcjmtdBtCjY94Wwi0/XoGolBd7ek6Q36o5TKVvfzWkhYDss5
4DWL1EMZcGcQkp2NZ7v6HI8nwccfbwRzpuocSR8fujOhNkwkoD1e1WEvIWTXwpI9NkJwbMPM1AIV
NysxEHGqubbY5793AzY8cLM9SRy8dVdXSa8aWRU5XrVQXAhAUdxvuCghvROAY5eBQd/kFII9X9Rr
8j3pE59n49G/bu7pqk3WU1eUzyFhOKb5ckhAnEXZOiHYV5LxrRSjmtinyyIbZuF4pKJt3HyIK3k1
HCJNr1qxfhLGZjX4XM7QDb9a+kprTlIfIZhVfTJSf8zkr2FKpHm7LRiYpulhATz5H1kgCsfJEBca
WU5k9rlZMRwpc9BziGKEeihkSGz6RiFaKnif3iK7UPwiuJcaE6j2fJACiN4f+eYphhLXQqSY7WjZ
FkqwBrWrAJ6zR6q0QcP1WrQbu1dZyYKkwhlHisTHQyqjp2eoFY8FBWUoJaQQd834VKXG4elSWZ19
kwxUmLBsSgU/OIdpkqenKecpMYpuBgY6nmovE4gA9DUU4QEEpYBAWoDAsny3Q5uin01VR9Ua8Zpj
L4z2Qom+Eb36tEHjBsM5TLPjSnBeF3aJIrhHOKWEO7IpHBgOfCy5EzHZqa+3nHrrH6/qqxMtEoWe
E6EgsVjQFbSEB0E/MZUsltxk4FsDx9rzpfobOz17b2cC6C/2K8c0xeoiJpuZFBrTMlUHmKs61WBo
BKBBw838Jiel6V2KN2B8qdn8vfb1yKr6LEZ5NKeRQWnw5iANJ/dKzUrdJIcpl8LFScDfrKjzUhgd
oOleY3JxwRPTHJnDgG5llRAT6Do3nRltN8+cCWbbSGP3c/+uc5tLYCjmjoZxlOxura1nP/X5z0vp
Lusv1CXY8giMvpSGBW9B95GmsgxgR0xn1M4RWal7hZ+6j/rKH03tM/tpRz/qm5Qwq5GminIN8wQz
KdeEOAYMg5I7QfAzLGAKDszceNHYhVoQrOlX0bOiptKgcjI8YhsmscBCS3L1p63ipqa92IFVRRMa
QImDOMLwHGPIT+cvZZ9QJWZIc/mOrYtNZ8nxxlUB5nQgEQzlFRj1BHXs0qQ/iVuqExFPyJ9ZiHSY
YNz0MdV4WrbS7laTPvDYuokG5KJ2Pil+ECOXCfKNIC9ObQ5g4cE48W3TbC0suY4eozdjgzwiPfRD
fukYrAd/UB1+T9j+ry8iOQn0C3fUDNSG6kP7vFBBqAy8EFaTaxX7mWPRf8ihxM3NP1R2E4Vhy3yr
MjnJt7oUB2WCrUSj4XntPBvG9+BIAaer9YiQ4A9WLh8bwzn9x/7rrGNPTlKSUJYkqXwI8Gr1nOjt
tIJiHWJ+hnGp+4mBA5oIi+yuuD2IWrUN7Pxe/38F3PRmmxiIwWoZ85e3KPtiSeczQN9bCyAiy5Dy
Mx78KyIgcv9gv8Uzz8hkfx81MpTGUcJySuTPhQbvuOce7sjqibtQW1da8zmJ/WTwoS0B0EbnkGin
al+jTZMSP+tCwIDSv13mHDrfPQ6d6s9p1qxOcA6dAG1YnQqiMFdC0Ois3NUI8c21EN9RPPfuUJGm
ukt1hOGvc5NoUMjgzl4qRFLQD6heXaCjbrFTrlHxSoOG2IJfWbZTQNHXHtqoNMWMGuBd/NnBTbMN
BmGMagJsZhNeXyfdVXPffkZeSZSslu5ofjIOhfitL+s7j3kRvme3muw2pjQskjOvkQE4PpP6UUkU
py05xpi3/mPESKWWaFUtk3HWcYHgO4ij9fCItgfROWPRwqkymYjxaKMpWU8WOzH0EC3Q1Xi3ekkm
jopB9mnwWRX4snJOmdAYPwLfk7tH9hUvGjSEGYzksJezjZ5cvhyUqAg6HLvPNfqLkb6BzqN/LTZZ
nvjI7+g+v2arHPbOZFIsmvtIctvbC3vK/tjwEgv+ufZLbtkrzpioEQCJs4MQuxVwgImDD8zkaLjP
ihRLTkpqv81+KQOEVqjY70KqDWByJjT53qmSrAe1z2bezfreIXX4ss5hXAKFHMVuG1MVKWUtkNJv
k9TKJlATs+B9Pr3r1bSXUBYlLMzt5gwAoKFj6Fb443tBToss77R08PjuojxH9kEkcnhVUAZeJhXe
Gs4t/bjRkdd5C5nK7P1Hv7g+TZIpw5v+3i4dKPUUcxA1wPV4Yj9SzFHv158Hz5bqS8C+PYD+6SMZ
noXIp4BgOcaiVWFvNuW+DqqvvIEDyVmeirK1XqTK/oa5/XEFnjVm5bVUM3a05qMGPWFu3MhE0gHG
vo7CzD6v1sEeDZUFAE9wk+B9uFNVQaw37exXC2/+VeIk8YfByi4DAyy3HQl7skgC34RGi7l37rIE
VIGxQCS39spdEdJEQ80oolIK9D2U4jhdlgrEWQXwNWxUZjSo0LfHBbGufk4U2FyrNtHlY/FnEobg
LH1MmYlNvlLY/0LlfywzcMiVbShQw/hvTIB3GvJrtYfvnY8xCRyaEvdYc2peC9pQ0pSXaRHdnll9
cOQjhD0YY7Qeapu4SRpquK6oMNZ8DaIs6Xv+uu7HGyYAUiBils0Xw4m8+V4XnKizwP/Xgj3as2Xz
S5wmwUjpWe+DPLP+P7ZVeSfTUGrx/TikoeM9npwGGvZG/U7XhLMqKe8kSkqWdKR95R33ciCH7mjI
iyZasm+C4vFMX2TPhOYt+G6MvLE3gS0ucDKq7pMZ/CPZIV6tdJ9JSncitiuFNRPpHKUfd8TNst7T
AiWZZoowwQYLv/yb3Wbwm1mC6C73zXrMxI400MGXZTj+cQbjBfasRoD4CrJyJxlSkEnF451zsKHy
3hByR/8Qk0TnT05ytsrx0Th+Y36FkHXTylr+9Yws5dUxUTWyC6/sBPFcGQ3pcLVuZN1z57JzZcYS
Q4xjBPIR7Rio04MUjRgxFUg5jcHG0a0zfntTJ3iPcyW511EfxKdzexwwb4vjbPnImDxbdduqqpQJ
8J+dFVZiFDe3XgHA3Qc4bi4ORhpDUTIchEhGLs7yBUL5f0W5C9nXLUCso2sZ08/3qkejzppkfK4/
PG/Wx2MXUTdfgGIu/WYhDohtdnAK7J4KbRrAw8Az9TNnCBWRVZEd06Q+Y+g4RH5DS7VUlurUbbDh
iUdmnq4kgCXNt2OIha+1p2U+qQxUm7V+6XE8/WLua7/EepDgYNc+StKXvlQp2479jnA7o20qsZL5
LRijkRiItI19UZH9G79EnpjG4LEhNQ3Zh3lWetM56GvsiY7B1E0PRN/P865j2Dr5JzNc22nhI8Jx
dh6q53yhub72xcLaUrtaoUjctszQ8D2H0qI/7nQgQsfl867cqOB2DvIIPKMWldKpNGAC+/KLOhej
X8OQwwD+iB4p1Oyx25v9WEfqwNCzPgPWP8VrjKw41TLQN86BjXQIr+muups+s60ztkBBQISrz6c/
zDzsLj7LjQCKvRh+efJ1tMSCz086y+PfD2h8tCS2F65KOx7HBsM5IYMM/6qwFOCBRycyFDhjZkYL
rXWpYwtdCzBbTvDY2MgSIkC5ZUeioR14e9ShDXJ7OXt5Fu6aAqRbTfpJlFI2oUekqMRUGhmGAqrg
yFPcK+KIKjNVeXdf4tYdIOc4OkD47OyigI6sZkvDJSbRF7HrREInRLGte1eau06gr4haXM0eYF75
sLbNs0L6KT77/LUSKEf3low4OcbHnFyUhuG7UkOo7L+SpChOF/icsKaJcIb0o7Z0L4OSL3LSiZhp
v/u0MGHDKkIYqBm2Vs/WRWhG0J9g2bdqxk6qTQePrbr8YNa4eU2iD4AFYZ4Fk/2qkaxXJXN7tFm7
nfGnyaUqaEkTb6KBA1xZM8UKaM+VroRgZ1X8h5iF5bvOXTaJ4JpzSkqsGgWb5uHXYUpBBb3twe6k
1XmhUb1V/0y4qn5brCOKnwraaRuOQWd46S5r/7KZ3mptzAeHJmhUkl1ENYvx1PLVGRIQaeGGjp1L
sLsDNULkhzct7DARmyvjoYbflayyv/f5K608u8GxkF51akGBG40NdyW2mKrexNUvwhZ7mQFvV7Cn
q2xn23cHVGIk70Ob2Z0HU9QPEqgre5NqU44LOkUrF1NkA0dEkhC+fepAV7KIHv3xAtnE0behv6mD
4cfG17o88fnnJPkN4PSHcS6rfoSYLzRU9DmIdADod+HcR52pNXSkDcSuRQUvZnD2dt62Wh4xBVmz
gQLVvil+bsXLssoyzCSmHv8WbhE0NLZZCWTz1M7872wpYYdu2NY7+Wpn1PrsQ/UpZFXUbjOwR/AX
BMFEKp9MJvorCKHFCtI14Hc8SvhNT31+tWWEAjyyDZzLEsRMPcEgO0o7WIdlrPnELQeUv4ItEmsO
4m5YwKn9RC3m1Gtz1UxBkcllHzb3jr5kw3+igrOC56E5oiunTvbKfOXKVE6H3lMCmZLygqXyfbMg
MKRSRiKWzH1DL7ajdYfy2M7jepXeN00bm4Jj6QGQBXbqtes3kKpAHmlPgtlf0GoeG8sT7c60zUy6
MdnulT3CVi2/uln8Db5eZtaVEW4ahRwl8ACgwwJiXpmn7pdI6V3lpf6PnikJW03UxG4ikN5wr3b6
ZAeIkmRvYxGQoaGb1OQ21bzQIvFaHuMYsvMsqTXs3ctOum3YUs8mUQG7/96/u27M8i+RYWMDAkk7
BIDxLEk29BKgXc0weNRsxg8hRITbpgxUYhGnnTuHURQ/P6HgzO7amkOtMPQeMrPDXLs8vFTVtkAg
jFAM4UN2XUNyYw5lzpgVO3ix1kuoziEgHUlcV9MrUtxX7826Ys5jfTGWhnukWhnQEF/nAW3EqSfb
a4R1K0I2fCFT7qJGVZp4qeo4dDc3Qu1cpvg599KgyQUkaSDbHljbb0B4kPsawrNwBvFFMNnSZ8Wv
1XNL/vqpVB/+7o9kM1PuP+9bGMHDPI2NgwjzQ17NG/vj93UZgwMMK6jANv7+SWaZcxVPFFVqg4om
kCfp0Sd/6zA65nZRzucCZ9gfOCwn4OkMO1ke6sP0AOWJNsdYd6HCetRdPSh2m/wVfWczQC6mAWhZ
vxNbyLOLKen96Rx7069MZqIArFKSMicNpDXlCUcZlkxiB4CjfIGAXj8GOUQUr5wNNMIaXmEoEIZW
xzcRw3FgReI/chMz/rPCcuQG+032v/qjyC/1bUY54jw0aFnuzPXEnqG9DkBYOVvImmj2ZknfjbZA
xrAOy63gbVVnhDSSHTPeohqnwumlQB1SW/sdUw6gWq8VvcoExVP0JXUdbi/trUlfn2AkNIODXf02
gccAXFoZVaHKCJE18n0gidlaSNNsN/9goJZu11AmWCOIUklYmEJ6WUVwwxmEyNAknWeyjzDngNQ2
IQC/tlEbU5dQBpbPZkjQzYBteyA0r0t9qHyaSzO0ZV7M80X1Sh4g4I7BQCLLrMQvvyLGw5GtzOtJ
WkEGh0qmyPkINDpi5YKSizhQpC5aKYIDZ/TkuslLlVy/gtSPEA+pdkXKhps+3KW0bUs+tPb3bPhf
7lDtza48p0Hxphl5wFSKyxNhBcTkg1XKU8gO9cZyDGl14KVQ/7oigv6/o5cgTc1ips2Ks1z1TCgI
XIn8ev6qxPnRntf1dS9ilrIurbBCYXMUDucgYaIE9lrz2V65A8A/jRP/WeM6bCYH2Uf30rpfLE2F
VAcAG/T4s4mLK3N3xpHk/xoybiEpP88jBTDZu0PfwaOvuWF9H9pAz0Md6ZKvgLTtoMVA3m3goPO/
ObrkrhWRGNW+Cc09E7Mu9zxVkzGWvyny7xfro7gF53wWbThtvm4Qiyx+OdQuoFf7IoGgNYt6zT+Q
+aGJC3bHM7h9f+IS7pQuQGXww0jWNZUfZO+gq5NkQXGiPsFBX+eMjcAs7A0QdyfiIyIsL/ztva6i
nRclLG/73H/eLmhff29eeBaSPohaK277KdB7I4MwsOC7JQ0G8BYLuB1soJ4OfxUqBFu4WaKC4w7H
cGNc2xslRN87PD4NZKzj72jq4kPBNsNvYk70z4Ru4/X2qYaiOC9KD90ok6Hzn83wsn1ltfykUaTD
YzKHgRJnRC0c2UYLX6p/eoXlB/PmS4gMBXvbfNEZzq0YwS3FmQYjNW3UtOsXolLDa1dmkcNrd1cB
zmupCtcIsnAIKEEJNpgCe0FIMGckEauEnr5CpIq/jQkOcryKbnWLemg8z2aTofMuHw5SRiScGa/S
Wg0m3+HbeqdtfF6/cwkk7hxQ4pP0dxTHvLqpkTnJbT/56HfGFKT031E3C28BoQVQg2DIntezTwwi
anybZaEbrxs69kZdaP/qDlwFDn/SkUsdqdeKqy0dyh3LhNo6/tgcyAhXxXF+L/V0mGndioQk0uDL
rQA6FSAZdo1CoXQajSpAgfnRYtwuoJf3kNkqBSYzx1ki/+v7WEru7ZGRyC/jxgBnPQtngBUgpCNv
K3kOuZfIXf4tvGgjMGFoIsLQ9etIk+jpMtlfJJ+UTquJxj2I9qkM1Gqu1OmW4MP6D3A1OKnPt47Q
Bj5q2PHYxG6KYiPiH47CXEbGXU0T1LMcd4Y+7Z4LLG3wWky47zIqwYLRPPRVt7fg0IzBWEpv8l33
TXqxadL6HRfu+UE4cRinFjvkZBsD56Pimtztz5HwdUGr7jaxgtXF4zujDovg7TuAo0y00MVFffnl
6J22/uDNUR3emu0QElJtwAnE9KVqrdLtRiSVKGR/+QjqNqjk0bCHo9Ffug+Z3JPqHs7ulQiEEj0q
XVVoZ608hZ740EeuUQVVbhxlX2hc4iUioRsfY1EL2xzXGYUKFk1eTDmMSjUB0RPTgcaiUp1cs+1F
AOO+2N9jT8R6tnm+ayggBljTuIp6tUlmD234ULznWNGADwnPcVa2XtVw6hi20A0sKI0pAaOih0EW
SDs/Hz4mXoMWmDU/2Y1dOCJJZYP1F0leHecpezD2b8Lbi406IzMnDYxOs/XC2yAzrzqojAxMHHhg
2oX+3R77eCSjiXbKplmUqcAXMwPQcSagYKx90qGK0q8C4blzA842LSyS3uM/3OO2/OobrztTI4R4
6dGrUWOQf+DGuO4pjlpBHoSWP9j6RRuSWWqYyyIRLrjYPZUD/h47QBBKpGZm1Ku4PRyvdQ6JZb7J
VLYj+mDWEH/DTwK6TYyEgwNCT7zZwwAKAtnE6IbO0UbQFDcspDoFhjadbAxJg9qawPwlPp9FS540
k2gQSREqdLjnq4YIhqsUMUX1JBw0q6CjFLu594+e8gUO7T2xIgYGvTaFh/AAes1l8RXoJF4fS+L3
xDyf1CbxKP/bUTPa4dsbAgzZqNP4nlR3QLDhw9Jg/cQkFhECh6btwJFYD7S8G79DHIAoVIC5YHVh
QMzp/zkqt7pQhIlY/2cme6Lc5/kWMwJzajYTmkRH1rqXT2jBv7YJEyVkqlrrFRi6P26NGWgADKJb
rgc6f7b96Nqr1w9anjtAuNHCzod6Z0Ieo7h4Isc56ekUHsQM6pmrIArRn9O64nw1l6DhSwgfDz/i
zZB4inAv36jX0bl4ZMq6rHz77ADjP6yE9+5SiSKdacXt+DCMGrX22PIrQEwfNp7Wu4ZOiJiYUZ0l
3ppTlmJUVVgvCAB/ROTTQSjikviuhe/IFUBAVmIsXWDZJa3+m8+UHY5soHiXf/6zDKTIzeyelXPW
ORfw8ClEgIEznfEkmBzwxNxwFoRaV0yC0AuGa4fRkQRwSVfIk9nKZD55ZczjBQq/1PqyJTrvMf5N
SCBxZP+SBvmFXm9H4GMmKm6+QaGIMCJjCj48XrIiDQ2Fdi0LUNSZA89mBZmcMhFQqSQUfGPF3SP4
oaXugDKWDI5WIWMQYBcUwnsy0IthQHoh7rnt9MtkFBrElbOx8Og8uXbpRjFjqRXEV6zobBeh5JMt
b53m0NUMPUM94W8TPs9kKid7Jbn8RW+30v/Xi/h58IfmklGSbaSt1xKaHDbgurOX3wIZNLVWLGiE
bRZthfMnnc5oqr+1jvcKFHGSowaLGKkmVSfS/+lhY6lzWRiCm9kL3OBC4HL6No8VlalGPG9nf3Hr
0OdFXOMLw5BDVLKiwI2hb41WUQqgROzRY6q3CiYbl+LenBOzr+5l7oS3wCa19gxOqc3C60YWOI1M
vyU67HItqUpcP9imIAUHWSPhInzn7D8TOO/Q0EYr5g7p50hHr4LYxlDiBuiUGSKZagPGTlLC6BVC
PsiXmIWMou28KjLsQU3MhI63kxBXe7MkHycabCC/y/Bz5gHKSosGuVpGJ/Sb7akE7kv62Y88EiSH
2oc8Xpm+hyS2mjAXnI1lFSVs2CDg4TR0IYyOeX5qYhCj0Bn1l3lLM2GVpkV7HMxzox4CgxVnGM/Y
b4XT3DovbPSdQd6GVtppYQ1yH8l3Jo9GsN5kV4RPDPCdwWECFTpBHu8YDjBYxdOpBqZoLmzvlfzT
8YHzuzW8+y+KXarefL0lJ1llk+NWEiHgl38zCRpmwccOGQKulpKfbwyZ4O4+U9m9bsCB0tqt/Ovp
GUnA18IM26EBmtcTZPD4xNvLQVzoW4SChTdyiFz967SsHCsifIyxdxza2cJ+WYRoVu8NuCvn0VNk
2qfZwkSQ3VHrJTVgcag7Jnm6zwREEbzadvPsy7wjR2qHAxy2H4cB/dOjzZ3WwWhb9vQW1R9VuOji
IscIb445JYcLprUknpK6MMK87LEHUVUnLAe7OOB8/KUSZAtR/YuKW7RsXuY/hYECBOjH9yKqcoIo
wWtXthPuDG0uo48MbisBrnZShI0VK/sv/n7zj7P3CORYqNlC2n6ttjjdYKcuixbUimoeI63kJ3Wr
MUR5qddYk6MyzWjpWZIcaTgxNh7Tsj5dh1NZFb3vYhfLZIP0H2qu1BNQgEINZ9LzQG1OWo0sNDQE
4lRfdbxe7XxwuE/I0Fe18PvpMB+lzoyU/O1iII5yCp01f4YL9N6bDV3wzlgRDOe/uoABXgJVehVP
43YGHSMzIKM21WRSEGwL9dfo7rUMo+TZ3ugSNLO/cSLoJiQVARvcphObroSEL0qcQILSLKlbv2rG
IYqjIHmLUxddO0XsIJZN7xd95zFX84h/hI0c0Z8xhP/h9UyBUYIw/6qG4KCRcIBZcKg7dUmLM7Ut
R0UALAGLubM/RFofbnfaiD73gM8MiApd8OHZirOa/3ZDRhGgYwGVSohJXJVlvq+l3+xUHpImDvA/
zHmzeTHwlL6rcyhdRVnI0OMIXe92880e1ItClcghByJxgWoviAKeo0DBQgqXDayTsYePOTkZLKi7
0glaTWFdZSDB3SgZSKhuvOW3mcAlhbDyCP/ofmLwIkFYkgWCDvWDmPFyf49e0uDarYytaEXCfW8L
wNnY6bGJ/8wlltT50aSVoZCbKuZ2yokE4XJmz4h+UH9qiaW+6aS2HocZiXt2GpOF7xSvL1ZZoibg
mv9wHng1SPYKFzRNQqunRdtFzlgSAj0eiFtbk6M4yu9vw5ioRdbAfZXdQn1MvIcNspLBYC1xqB2n
npv2ie8Z1uI1NjUmyfp4N6sNL8DusH/DCuKP9L3a6neTAxUfow3FN+TUNtH1HqbzqZs/P3XpUGI5
orhUEkLX3VWMhNmFEZcmJA17yiGI9oBit/clYIlCf2yK/ZRvovpXj1w+6ddNGk9LYjMWeh2zVdGC
mCXGKGArZfxQURQwh86PnXjczw/WXIMJ5b08NVDFJnyfRLNPSFA2PRa11zxDKlqvGdDyiKy8rRNc
jAkppC/rvC2ojDw5F50UAn5T3iY/jzjusDNWIxq5IDGcsTvomK7S5KioW1mOragdVQELY+hdf0yM
gp6v7uz2vZIDqHhkUsQsyWfLP1TXMi1XD9YIajLb44M3+KkNkGS8LCjjPTW9JBLyjGAJVh5BoD6B
9DWk50658UcGhoP1QGiqw5BfT0Ksmya+YoAw/jY9WHMtqSLWcOSMbVIX7D7XdwqZuy8Gkd1EOaTx
07RtGV7+EQMUp3AxZvLpUn4SOqmWVb1fViGp+ExKjOogciIyaRxTuvpthcXzO83QAwAxb2IKKjFC
pGI6ng8cu2sYUCK8t8cmUnlhXT3c3jd4+41kWXS9IOosIMkwgo263s5tU5LFERP/IJ4uWqsjVbYe
g/FFlSOVOg574sbN8kigW2LIWvRT+G4GuhL99XOkW1ixWQ/y+5xAEQ7lRgoITmNimDgO+GaoT+cm
D0MPGw/su1+LnesH7Qxwe4ogKuDTw+VcAS6+dVkQZR/1TROGCW/jCMXH1bOR8NMTVdmVGNKgmKQL
opfSaTQ37fRQKbhggCVSpNmaVc3glg9DxFoQASRIj090IcOhEnb7jOVnvq+hTo8T7Lrbpvw+R0sg
7qqbzqpqgCxxkX6B7564VzpJqFQvFotbwMg5bRKMu6l6oy7GDvN3ECWxMR2WFmsdfYeDMkQVRzjf
gwjx1T2Owe4Zf6HYJ6L+tOvM12fx//Syod7ENkAIZdKLEk1BrzDEsLsk1BtaWmZRU0qx0Y+RY6s6
bba/It/0T6GX39UniSLJPlyc7q9uOMrQURzgnJHrVAmUZNK4wQ3qoz4qwFcs5bvvmeSA3oTq3pVE
gavdPCdO7ShXksyQH5tK6xGU3F8esAArBwqe9wrVWu2lkO0uyrQJ3xU26Vn36yFReSiR6xToBpwZ
RUSGw6p1PgII9rTX/W6eFRhbSpj51F7ZmVqcrlnerZcN7aiXO81WlYiCAbBQIlExhvoOLiTxXYfw
m9G4fylrjRL/7FWNYlxjCWC6nR7Iv/HoGyTRGj+cx8dbkCYp2xv7kEuDoj6hdVaqOJGBHKCb+LKp
NzHXazF/itqAvaq5Cmcn5mTg2WnYyhYnQVqbG5qLbA7ffVpseIwhXESSOZSAOKrvIxyF/0zzxtJF
Ujehb65HFa7RZmuGyoOgTWmg9hRU1Xb4AvlBWkSRSMw2HKfF7wSB6bHb7cRAAW49uHyzfLa2UMZ8
NbKK+cisXCt6OPx/xv71ZQkgPowIeF0hEWZbPfjKAWGaMuG/ThBAv+SfODm5/2DRhvsfbnDrVRj4
/2IeRcRwheFZRKtmx4+Xm4wd+cXVN6qBzWZxU4AeoEIhTks9VN/etczGzVF7eTCJnYkKpQn7ULE+
Um/pKqSYSJFUPLMG3urHw3BB9zx7/9qbQYGp3zB03SpL4xDvWm07nv6HW+swibTqhM4/mPU2Ai/1
iteotxuWGF3IreNPAGhhDxOpVpZaKgGPEOPYuYDgQcTRJqe6qvC6yK6s2TNbzOBs/StBNyIVLacG
vcd1Vxt/w3p5k8Ne25gOrPfKCVxR7p7FlTO4FbG93So0oEWh2iwnHKPJ+M6QKbYQsRYxng0fsZ8E
/7aFqS/DJHFN13du/xapAoSg0TwzabEIa7hgMkMKR9L9qXJf21NVsfgXszVDlTPnzvFvCqYAEurJ
exkbrdbPVhR+jaAPDK3BM6EjHjcGDyrn+BCUdX1AZ1Z1+ROv14am7W1NgntnBA8WA/J9lPhaaneh
Caqn4YK7OviHh/kfHIZa6TAtw4NdlThuqi+72LgyjplQHA31lsZOE/g+LitPM2t+TR4MaGlcaUKe
v58vdUlGMmziH7Dd01Znc0kjo7HQRpJP+gaj1t7dTrk1Z+ebhmFXngCZt7uLTwL6f5LMXQKBjy1t
tGDdmeD0mRc2DH3+Khe9T6wC1gwbrie2WZZbsIsGeKGCcJq9Kvfyd8Qvohd24UQk4JSGflR85oLy
JDxb+EL4mH4+cOg2yy5+DILfZQTM7ap5sb3ZvAPooF3fbxHyHUrGHvZmQTSKSoDA5pTZHhX/Aog3
kxMOtUPktyOY5rboQrwbP2HPsRSQjK+AZWs3Xfc+mfNAoP8ZEL7BmlL8MqVNSFNuQVIdqAou8l1w
kc04+mbUnZ6iVavaxQFH14K0LMg/aiZTEovt6RSATBsmhcjxFV+XOktQpLxS5E+pkJSaRjIuH9hM
Fe6RRpr7Mt5C/YIx5VbW9ZNiWyY8+6mwiKaFbcCCnNtznvTie38iY6e6kejesf14LWemdV4hC8DL
eKBW0hZ12IO4DV9FLiDc5+KsexW2f0CASLoXUooPDW9zMilBotx5GEmr5wbqSrmm3Cm0BcH2vLCh
ynpQr/xQlDYEy0zb1hdAYukmhsnt5ztMKW5jmAGwTWJkHYG2dBNmqWQD870iijA4xDQTb+jjuPGC
lYAmFiVjmvZbE/11uykhKHls/jYYK3vJ1odhaifE4ngewpnfX7ZGRAJFmpd1DWfBTpxlt0lHLY/1
efl842E5SlKOo8MSY2mnRmP2f8ZuvgWi8vlN2EufBUCNSSWdSUaEkOR71OQ0LeXGdMEO6S6cFhou
o9figCtZ+QvT/wHP89gJ5E8oY9xYxKjvZOmaHTcubZy3yYysQmwGNRsYIDTYpFpSE3Atr/K/z1Ky
zggGx+68LxSu6AhJhzTHA+kM0cKxPUvQMPW4ubTBGiCCUAsHoTBMwYO8niNvFm8MasHYXRVaOS8j
WCpx1qZOvyzOnyZNN3c7uJbf6zDxXxGOlsqPFCnUoXyt2NlwDwdui+xWQoLhPgG+rwLB38UZKBq8
xed8Sj3NXibu9XIZ2NldjOjDRMOqNFNJzHG+IvBlZiekMZF7wusTPIbCU+XeOn8kgzwJYyE2XF54
laexGZkPlRBDIWhW5F4s8UA78H5/6YlUbD6m6hZxRGM3w4VBn2MhGjeJVzDd4owVBlr4TjV8OOCY
bP0zO/CZ7hxcM2cbZKoRyjXhRh/tpUG39bcvC9K0HAlLFvXVzhYfq5U7f6kvpWKWxkvvCnhY+mwp
CpytH1ahNMovqPaHDlaz3OmffbRz7dQYfEXND09Aw8QZ160HC22cWyts1GKaPJsqKYfHyqaF1DWM
SI+/ZYM/h0U4yhshY8GN7VyoubQthpoyN1J7XrKdUCujsSjRn58zz3TMJqMGdtcbCfs645SszRbG
eZ4X7+jkOoBKPaebDBo3GrqvOgX6PJG0Y5+r9xXDMCBlzsMLjjmX2lIgC7Xb1Ss+/I36h53m8WRK
ArSTDf1WT5iPbVNnvtR5Pk1Ey+yKq/WvgzCOCCW54pB5YJ+dK1cIsP/K1SKxvc07mIDjJ0EG9KXB
OXIVVcpDuxmPS0BiUV+C/lw4u1ah5HWhSxk8gg==
`pragma protect end_protected

