`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
a0qszlI+O/DtVIpvDOwOJ4UzEVRmwnhjgA++M0sJPiU3vTUdijb9uKX7FYSqH/VZTWIrdG7rjK8/
aQjel2mjF210Dsy7uWw+K1UGjDsGQdc+LczxDaN7ShHcmiRWVz3cxHHoDPsbukYe1ytb3UKFlwMC
n1VGGF4jVyVrb1PaNrkkAvNGEfo1+d3ItaiTEMu9kfQneFPZ0g5Y2FAO0bzqDlKbIzAgr5Uv7WKp
+0VrBr/g3yyRK+NYNmNq+2RSSScCdqkfNAUNPbsp6DXWjHTj7DrEl/QYzo3h800Llij5b3pAS6Qs
jP106myo1V+PTfB2JtjBXBVKci0WVMV4HH7FiQ==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
xuUMvAQ45A1fDht7y7COpTXLO1RSkO/CSPUpuHt2EsJCDV1Sm0cy3DvcUvxbfAfKv/k4z/ncV1CM
ApFWg/My9sU06qyMjEmRSX83Me2cLDgtz/WKknXgDD78fr8tqKpd/3q5vMD0rFxMya6r4Glqka9v
3kU4J8Cw+UBfcVMMYaQtxy+qD1ZkrQlV5Rvl2tOPB88DesIKsaCMoE6i7DVTcYIz2ohnK/FN+TSK
w5F9u4CiS9y/Qw5n1EFHsLRgo9OaVoOTgvU9GjccrVrD3jmrWAozRryLhdmhRwbA1rw0/SryS82L
Qf0KZHZBcg4Zqq13QhjNZJmmlcdBIJeJXCqg4QAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
oQcKNx8TtFBUWxvcIhKWUGrkwIf0l+I6e+Mffmwt1OslCfKGgfF8Rkn7dqCjTPgr+/bcFv25+57g
1wW1FM0oaA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
iVnVBMoHtiJcq5nXtIappPv4Efedx2vJTwZkxKID9aYUptwnG9Cx7ILYxInsVYxcrY7MDqsa+b9X
31xyG0N8vX2esSqwuGOra8cEyu7jgW/bY1mR41DMuRdoq2f2rq9VD+F3dWzpTBrdGgIEhDGQ8dLD
GEF/5yo+kaKbHaGioGe9A8XW0ZLU3wnGAVNu6C+b56fvYmNGNCJzpViixxJloN5NWv63qtI//YFP
o4B9Qk6V2daGQZnOZYmDOagUWg0R1z6oVVkr+FpvdvrouePIIsYRV5KiZChiP+iu5zqWEoJ6v1y7
68F2wGBucnvSD6QkL3TOqMagSTlXdagmi8I4Ow==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
B/pWKO27dLHuoSKpZ1V1kqOra1plkeHHcuikvgPZF+GXx/GDHIwWRKz4v2IgIBCZrQnJIttu5+Jb
ms73K6c1RYRKHzWfj9FlfFUEbLW9W9bwMLKCm0QkVtMtmOVT5icl6BtJwNYY9KBhFFRWfmw7Z77z
i/t4s7gWQzbvjmzGbLLtZwKBL+9ZFkNx2zh7ybqDVvv7ZaTls0D2t9U5NYj6ALjYdv8YRnroZWko
UhF+KOM69ItznZnZ50B1qcMlTolGdYVfo6CFO2UjhRiPttqDq6iEfgbIRtRNbTi7Vj/FNJeBki3d
w7zeC1EGDmdRVNYuqcY0sxPTavx+sX5ZfPCUyQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
qbQJrcn/N7D9t5fBiOfgXcEXk4WzQUfvveRvyICvtyk90V3kaGRO6MThAr3mSqvcS85ELFF0nKs7
ro0fgAJpuXbbhrcupfVuqdCYIG/KThMuJ1us+teMYXNkPpyKcre+TD4jSW9wfAeQQkW+z42FiHvQ
eU5wReogMWXE9iDJXmg=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AiTx4nCGd0GMk8Mn+/aEJwT6yKklrcYfvNVZ1wt9THylebRph5Mp7WeqtvcARmXu14EqpJ5aQ+Oq
b6kb4w1L1Jm23fwcDEukehlXuaWipnzZpE1iwWFR6YP+DLe3+QY/ZwA3nJyk/PsMeq3zf6W2l/FF
M/y4LkpAB5iLvDjD6U6yzokDwHoJBzrcnp0gHhInX+Qo7ttg41DlV72tQT6D1tNAlrlHqYEElyse
ZJptD0KHaUG6Z7FDDMMvoV89GK5eB5NCJ1gBIlWldbilA5++jmIesrnhS4QkbLjS3TIj5e4778qL
sjqGVQyAGHQoUzGWiaJmSvQco87d3fpBRjCpSQ==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
S7xqXcW4TrXiUqO2UlDsoVwmT4ye0heCq/C/CsjbdzCHt+xxHMpWhu1RjHgMO5KfsXyOxBu9txnp
uX6WBiB90DkLgmbYHAD6PMhEU6K/jMhe298AIjKeKt+DzDtQYdqo2uGHTygAqXbqW7KYPwZbAE4U
PSHI/rPlAWHnu8W187huP2EGcV61P6b8l4fSzOKhk71poZ4SswCa4pDsrghspvwg4mCufurB69CI
Irk6M75RP4uUSPv+KULzjR/kRhPv1dzNqTqwoJf+QBfv6yRB5vl0GjIkFYd5VeKHbHDeDJkD7Rk3
9cmpWzhQFqXOWaWa+eUgWDXwm/9c2/Bux8jk8Q==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
QMwU9bRZq22MA74cpW+n/QTf7arzUpxSRZFMpi12cpfkR1El+lTzr+0DBEEPgcenQgcHT1dxIbQh
xYFcPjbcSeF9BVVopfHMgesnMhqyVDtEMUDf5aCH/tkqVkjEvkiqxuGtZKnz61PHxCatXeelsSnt
zievHnEXAF23b12TMlA=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MdOzaEiZC3B32CXoThl5o+jOZ4XNcOrROGXtAk9Bvm7F5ixw1dZYp6V/IgUzu/YdNu4MAZGh3qXs
dzoNhBQkKKykSsO1JNwDeiOW6CFhugleitcfPFdynkeIDkoYgv7k3QlzI8kR5PYa/Y3Vo3yZJ7Ry
B4tZLpm0JvgiszFnHK5Njcm0OcaP38R+nU6YReS7pqbHhRhA4TXEqwFI06VFrO6/u9EvfSBNAAX1
OaYZPDQbv6SLEdJaZnQfgpVlcMJHox1Ifwzf6l+TqPDE3YT1UfGOrc49RqbwO0nBQwRvikJYwQvl
PMHZBPub514Z9w8Q9j0lHIummUKAVI2sZBOzaw==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`pragma protect data_block
OLKst3WQdS0v1DXqOEBqM43uSqt4O0olElbuVhv5gody3jT574Rgb6nTVw3QHZ0+6WqCxs6aHSol
NxGYmOO9O8mOMvyzo9dTPjcy/dCU8WPHPV02QvPvvS3DmVXtu6w+VuvE7/meHCBDRuUQqI3Cwm9E
H4B4m27Og9WaIjIXCUlAMviQnxfPvZ0t0GVEhxU83dbgCMMPd0lSkV1LlElbHIfIqhkKk9/75PbL
HHagB0P8MXDnNFUENZU5LJ1ecFrR8Vf0VmbsOhxZ35wwffzvaHHTdEXTmZ/Rx+6DETrbGC53lKeY
eceLIrSr1EIdxqT9Cxgc/ILYaJ/mim1lfKqQc73fNib+tnxe36JGNt2uUI3IeixQWWVNsrPkGyv0
dp2CosivlPQtwmfbwKq4IT2MIS2hrO93Z7aXArPvdGg/rLf3JCbk7CGUNf3ioqUmtHDUbbh/Z904
TxAedYvpl7XwdJIGuCdYir9S1GMUhsllSt2sqXxvDSC3lrFBAg37ON0gGCyy3okTiAFb/AuMOfT7
yizNQrDyAs9HqHHs8tG5ToOnK2ZTaqkzXq/4M31HUj23Z2ceHjRqsXt91qjrLtSCsHFLM7x3YK1v
rTpB3X39j9MZ0hvtZYLompsjIZNuM3YaBQ2nKiDaA63RY0B0snsn7vNEg7r7BQpz48SQin+RhO1P
xXaPFTBy/61rQeW+yaRK19PAsF5PgO1pkEw9ZRfQn4ZjauYXPok3lyK5/F6Sg0qg4e/zrNC66+9T
gASyqDIXcRN8b7TN/q2WUQLLAeaeIMWpC52XwRzxiAbtMKenBPjAM9//+gI42Pu6fnYa6E1ZZWLT
3/mIsQrZTzA39pwF7QauABliiYtBEjX7E10IJsEszZXWr9EMNIf+EXvDJwlFDU3jRsdneBFTd3QV
qQL+gJgqIy8R+niSEIMqGjGS9sqG5G4K30iPx4adQgAGx5Cn47yW5lZyPhGbByg7i6BEui4bkZ0p
whaQMd7PG6Vbi9IfbCSgR3/zPpyA9bqDXbgH30wIMHfnfu0o5y8Nu1VF2PSjl+rDefmZ2iHulTNr
pWk9X2G1tabGjaDXYsDfZPhZLJ+JwuDQ4EFrNaRmcv71Oj1hB0TnTjYmspvPO4Fnj9veefIw3ZWk
7OWk/eL+60Opc948yTV6QBKPpxiCV5KffZRds/WRONk53FIpOdh05WCO+7ngzzdfOY7Tm/99/42u
HpCTYcUsaSyRCqOWYtFcqsDp2qWSpL4CZlU5wDF6fHjC1yioOvwTIEwZQqEnW8rIYNKglDftnZOA
1XM/AxCw3o7BVtVAZOCt9OusegcKb8LRhyjsuB7M0/UUm+EqOMFD8huwAiPyCgTm/an1qHYLG9Wa
JLX34pU1fBlDd7wpTGwIvGN7xBpahkTiXShuAUX06yXTAJgPwcXr4qwOQxfTbRVSQSA4/xNdClRe
Pj+KfuyVzPgZZvpG/hVe4gwwoABPrWy/z5n3/lZRLS/fsY44ZdPU2+MAM9ktsTmyvsxELOPDYin8
+lJl733DeevRGLDlWuA2naxK1oS/eooHUrFJUi8KWQPZ6FIM/+snzv54O7x2zoDCx4kBa69eAzdz
LwF1h314BaVDFmXY14YAuATy3tENi8GRDh9lujBpaUldgtt9Py6VQxId+3Zwh7m0UPcPADMYrl/f
0RVzwlc+Up93NEzfwEXoGqLAsYNGdMKCNa6abg6eSc/r8xgnxK2ygXAQzrtbaenccxAFtNCCKOGb
AmhhK7dMGmUiCPA1DNTZ+GLmr8b4xSVMiaPVFFZQ7Nib3eOzhzrftfrqCjNiscgJox1iFFDLk/RD
9fw0Rs4gkCerHiBaKBvOqEpC8nQCn5f9xBMUHr5qGtaShTiNEJHFfl4YIJ6XtHd4ufysfslfKUEt
fiE6YWZgfLZoQoni+n/EURU947qrBpvcocIOyiD26b/HyAyXk4mtoGeIIs3agzd1bVAsTucb3wZw
KqSn6XHWWt0kygtUFiki0I0NRC2NEGIZnC1Pmrr0M8R7UmjVh0KjEkW77uywJ2U1z809yALeIkfW
Jfsqtf/O5bXANqiJZjP1wea72RY0L+2aOCEAmzyPKQstX/tsNRM+LFF2nj9Tf4SvS4GFflmJwoRQ
IdlFrCALS8iS7F2Wg3XlBXCV7ZI7l1VIJMy3lbgykKJebUN93SBhkZtoZVNeN/zTNwqxffYp6sWr
zPpp6sQqhF1sWv5duWJqtbTRsf25fPKF8TZQmK0Ig+uPoM6e55fziBnDkgGkNoH+lpZkqoihej0d
BolhxA6TvolAxzMRBXmnGjKXvcaIEU7lmYOeQYIqZ37+Ak//7CjIlvokaNewBhhc5vtMuyvACkE/
V2PSP+m8ATvOljFVc0v1RM6/ImPaT6681MucuZPGUAvwBVBGByd/U2EWNbMrYMzjhyswxB2lBER7
x6EGVkLKGFk7wSOaWeFpC1Jnrd1kX6EYCftyMKr0rp+bglkNfYIo9V9Vf33fZ5H6RXSD/cd2miDC
fY5fzcfw9r97XF4QgW0lCi6LZmCkHcZlvUJiMmfNmLAziUomJODIPhssPxndwnFUbkWkXGb9+mq0
D05WpEHGFz+2waGWWWL6ihimvKfRBiqmGq+zs65WVRR5Z8+oWNzAVF5AZYCuU+beepbsd7bi/kLf
l6xpFsCzaCzhWAd0smT/gWUrXkF7kDLsLBZoQ6ZESuDrX8Mds1BlAg0lUxqXbjpfsenUqmKOFkcD
bowIoD52OkEv+MV3Feclnhnh+MDLNOpMSGYBcQncSBJRXnNu8r+aF0GR5laEb8ixgoXTnAAM29pd
b3MdaxU4Wuwz1xgx5OHo6GsUYDCHNCwdoZzUvmcjjvHGiRQr2PE9yXca3llbmaPQ1YMEaGOmOf3j
luXGWgTXrXvqFN/gbTQvtIhvf9mK82h9op0u86h7VvRjHVWRM0dikexf0bgseUFgNvt2M8jAIbcb
y+DY9l7VZ5FCbVmQeijuvKIppktj4SiX46Q18uQ/3hZwhlRo/7SFsQq3JBcfV6MUderx5dsOd2yU
rRVwCwMT/aitiY9CBik5SYXRvbWl+nc2nraEMjMd/0SZKDusRgn4rrjk/PBovYeaR2J9xu83B5Lw
ILfCAcIYR8vxWnwi75P8751H0TewzNbLqm3wIr4gTwmhrFLTqnOYczZT9Tw5wZzVO/9wVh86alrP
aQwZQanfaIABreWFeYv2uZdsN0T3MNJYAOUryRhGN8QGHeqdEUjUF5m2fq3OZZbpHbnOFgEuiO2X
n+BxhE6pYgy3ii7HFepMD8ak9hd8u+UhJgK9/BNOPdau2uf5DXgHWzl2NjeI/XrHGKAyKdex/7XX
+RQUqywnezmjF27F9MGFqxKh5tGVOoxhiYiAAb4z5QsjqlQPV7ku2N0UTK+VxCapGJ220ei/ZbnI
NEU6kYOUePzOWxQSfolDvlCC2batcqaKODBoGlbxMIOzw29Q+y0ik7hm2nvOAZBjy9pl+IirZeHB
vawUQodSTyS415F8eRT+5It/rF06LUj6IELTEwENIzp/HpVqe2e/tfb2re+bvmETx6T6Low0ZNNR
osNca2FQpYM2InXfi0hm78P62KAcE+ULnqEvtR9TpKUroTfskMyLeL+vKA3YiZvfbik3LSfHSHOT
/XXW5kKjTzhnoJoyxeodFh90g4j4k+MNVQZZFkHAwa45bEIMYXv0Z5r7GG0NBaMETwHBK5+CM41R
LUS2hRrG8LG16+/FJy0c4vmHMUIXohRxxy4dcLtX1wko3u7wqV2GuqViWWO6sKK+sYCh0pPxePmY
WbZ3rQ3r190OQdN4BMIIztqVWuzwJ8wosWPeKyU6VjZ8XJKSSO9mM0LI8G917ay9iaSAl3YTtl5w
zrXdFeoxM3KUnYzhytxF97wxdEw7FHdaNOJ2HJXiIse7bgv4k1f0ZqAv1PX0VKBTQ9Iu8c2v0oyL
bheueKhY+ZRJczoeYNJR+L+vURx8QCNwqbT1tH/xR8IaQAC8xhhka8jkO/SZVNxBWrXJco9ugIvR
i5272pnUvV/cDPK8RrMOK3PhGmlUbPpUp+WYcULSAVDIJL7Qecwiqkn+ncQgy7BGhC1PSoynMxHW
rpONV8RfkAw1R/+6jFtZjyhrXuqKTMMdkEzhWd83KzRNssG8nhaCIXVu1GMauVqxzMCt43SeBVLd
lJrNBut06YiWmsQbbZVYkMi4XggJHKgN61LFHQQUYFKu
`pragma protect end_protected

