`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ehdMVNu3vuf4CFn6zvT5hrDLCEB0239WSkPOw7p2iKx3tWdFSTBQidPZVbZ5ZySUZmYIzxKAFSLx
x7FoPYsW2xWAiTi4VxW0r3P55dE313L1BhHCXiBQ4qLTxUhonBoZVXCyfMji/eZivxa3DAsMlLtG
ZNLnZnsRHS1meCRrR4aE1aFLrPkE8LPa8QtgfdYRzAAct41+14+mKcwQQoeits3ww69w2MHS2tza
NW+bgkrhPeb+rORPE5jA07eQJQseI1SWN0NI2FKa7V9HJfFuSFfNLgviuprj38w9lPzeldMCZX7w
/+Sef7vr9QoDomFMFGzzxdwZXjRXCQO00K4vNA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
bYmG/j0Vz0qxbkQRAcBA1p9TwMqcwsen3xRCaErkJmXArlRKWIxSyc+cp1iZwYBDQXOyj5O0i+Q0
1ZKdx57zr673hTURqZoz9Ts6FuEnhPruEnKn/ngBjc94xYxmmqOT9T2Nux7v0X5RUadNgQD55Ck5
o9CT1MVPP5lhiq0ZlWvjbx3y5aQVLyqfkX5bZ7lerCrIUCk4Oim+JeR1oinX3f+4B8jGVNkfnTZ5
fqJtheyrnvAYfwgLRFt/QYrOpSORkEppSEbhEPjhTbEfcM8c/smuVot/gzgT4FZU5D1f+82Oqlxs
X4gt2/FbVCs1Dz34h43BGWYzbjlcOww9qxewoQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
qBNrVXbrLGIwuvMu0m1OnFn2Q+e3Sv19X87Juspyx2KDHjSUNDWhyPQlcHAyba4yIGICMEdEvJMg
zIUzArKD/g==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
QoBTbh6d2G1AlCMXSDkoors8hpYdKKYlqAjfdm33x2VgilBCTVZ7sf9lOIRFAkyTCtV1rRX5CrFb
iKJ20IH0ltHB1OouwG89PWa0+RfDQxKLeT5s6uXKmLkQEu4eXWH65Zfy98t4JrbxRyVh9W9DJr5L
vmPCKyT9dyC6NTmnvnnSn821Cas5O4uI6ES8riO/zsmsAF/xQkyKJpEaInqJTZTOVdm/95B7tGvL
LWtotOtmCCFr4zYXDdYT4PdQ2mMY1XiXIVOAfrHECtU4JlBuBj9NUP1c66rlkGBp+EOvclGgpTFP
ajAUNV85Nj+DFKtLjsOuyDM50wQyDVLj1Omjfg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bu7bhcGcJAMUXYp1yXPU+V7yZZITMHlXIaJRtN+SB3J+s/aGYx6/TMng4nXWtj6daIf5sKU3kj/T
q5JVQ+/tbsM6YZcSjvIfCZc/hKoe6rKSqNAer6gpAjxh+sKYBQq8nEUP0pijn9Q0c6/1v87o/2XP
JlxIkZzPUdN0OSPnmPVVWoBq4ek7ZrfYwqFyYu6/afYjy3KR7eAdNzgWEZXuPu0IfA9y7TgTUTYy
5EfyqjRAoMYZe2EpA3YOCbTqo3yf0g7HfIc3jKUeQXKYaNDW3GscPIwY1wwVzZa1T7TTfsEAjosL
S9H57h2vPV9oXR6+9ctB8j1CfuFNX95fw8YYgg==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Hvov7LG4UgAau6P2mLIUON5Kv7hfXcnbx71VYOfp/D6yT+fSP44MecJk9pP7Hi/F1GaJ4LCgNOli
0HTopsX92QYdnwq6EPKnnyQNbTHsMN8ee58nn3Yaz/VWiJWYr0pm+KX0ky6nqHsqXMwBq9KHvdqz
DVf6hIjO/wi0W2c+pgE=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ddSeFV5NIKypKxkPzRYBNWK9AO0ygM1otZWtn1SIXFKolMPSiViDla5H0uxPk69LJXqDetKDujBG
g01FLbmcLQbZu5gj0Qj+xqngOipcI4VTXlESokfkcca1tC/DlRK/4dxEUHxF88AxDeVK5ghbFRV1
fSHmgXHKxnFQtnit6S83vrRWAaKSrLnRanzgpLXogfnVHkX/yRqXsumY6fhVDlux1N83PCG/tBFh
K644w1TKVGY/7YSvG80nVoyhRXbpQRJsvtZ8enhBZt0weGLpfUgBXczslmIMKPQXDczSbxhOGsni
5ZSnPQ9kO3hmhpsWMLdv9vG2Jl96VXgDeadGKA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KafrQPOaclQ45EUBbA0QW1t4DYuqbSwafRKnawyhYG2vj23v5aHYfoqIAah0DEPfEQGG8XOWBlPJ
9Gnv+7q3Jm+/VcFsyOajBxsh1lRtEGOo48qfIG64Autq/f4rLZOYaSO/B2/eQ9P/IicG1ZtX39u1
Qm2ZyvvSBIEE2NYf8UfrdBnuxNFeVT6656Day/26vCPHRSNNvlbCajEC318UF8EXrKjb110lGlj/
OX2zoV9XMwnQYe29rm2VizjKZJvgIJWjxVzm4vSglO8KYivzRhAYeERoSBForkWwBXd8CwwOeFzo
6G/5HEI3SmxzkPGkWJ+RcZE5npVpxeNjZpXqdw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
N1NVfv71Z/eQLtsU5jOZ/zJYbkpDDbKPDldsB5uNCXy/tvHTUPEh+5ulO7JcZn6Rmwq9sp3du3b/
MdtDA8dHi3tV/uhHdpvXN1iD340rjTZORPaypB1aAacS/LAW+6RkK4QQmEVCBiCkuYUOAPJEc3qt
aUq1zYmn5tED2rLmrag=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
P+0ACIXYteCOx/Lnae2cAFoKYvCHUBf52WRdOhtLw32scNTkZFzI2ernJx7xc2GExWp3aAwqmILm
bGc9AINbhdw0/G0ar4au93HM3M194fvldCAQCCK+6WeSU1zPYw1Thzf+9liC1xWPsb9fPjvdShBK
5uVRg5xrLU34KdHJKfsaqUexVXP/RDq+aFwQYaGZhzLaFg41VjrXq7GSmhseTApGS/zEAQQZd41V
78IMHxEG2wC0wrjYWkXB4flzYkhNiF6bDs0uUCg6M8CepoHgYhVMt3arbpyearJicJN7j7+aDryf
n3Huwc34aDxUoydSGViJmeYk9HVIhpICQE/nhA==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36992)
`pragma protect data_block
17vf296iqHM0YYbkCjtuHAiziiRxH+0gfjDBw9OHD+fr5hkG+bRE2hYwOVzVN4L/4itWVrUWG6vM
bu+Jzp0iNI79ieBI4MLHb8OcvKFeoosz205WL8YvgfOtal3c20g6/zDtjsCGar01dOnL/6b9NeDC
SujtlAFy930tI0npLWRMYUhBuaXHyIrXACeAFZzn+ZnhE9BSGm6S73RNF3MpjkVSbCY/56yiy+NT
X99m/FWNEG3LLRZxww9EQVGplseAnb2glbuuuH0PhgqQtPv1+1q6nf4RIo09IEFf60YF7xemoGSM
HRQQkhoV4SjBivOPzLZsMwUu0GPrs1pQHoUX3KcVcAPSqhKpBXwaFZAZJl4xUpB3UTsRmrcKXVBx
6AYj9v4kKrn6pG13AwvM3ieRgccRjFy2nu+LqcnT1DDSySKCJ/1+q/nuhBcnAVbSo9C6jgmG04tJ
jaElHlyL8qm/kz8XrXR1C7rlPViYc+aH7/9fdf14DO09ltR8VpIcWkHMhEcpOwdb0e4ee2l+npjE
lsIykk1UyVO2lY8ZwSN049nSqnjdnHNtATmTzwu7Nq/oehbzG5T+SWdEH08IXDBnnk0DKv79qoRp
+29f5gYQo2jJyCAL3ib0HrKPwydWRD41Ua0KHkxEgyIVS7LQJVhezcmYu90UOxyKinz2UNWRbxBQ
EXDTfoGQYmIRcdsqIR4MaV9Cb4fjvarTTuLpMPCPGtDStBH6QxvZOeH2gqSCkBL1cCeUz4w9v15O
APOXJkK4wjXmbqkgEFCSz/wzi8I5bxIDVWnAHyU3dAEFylybRNjOkUO7GBNL12ZX7kV9G/U0ZYsK
O4oY5pHfn3fJXxfK6HmvqajVD4EsJEjG8hr6dmx16FIQYmamNccXkNFDtzmAiaukUWiC2j6HrAwg
4FUpKjTEY5gOfPbbGYoImfStwBZIP0VdpGQxpkbCf/QMbF3U+O06ZvrsozsNNI8tS4y7KUS27z9D
IbOr9aKDJh7xlO3waAOvxS0Ai3mmnP3HIljtDalxPIC61r1S/kqgpesDxHyk6U8/UPzWUR26YauC
mHUa0iBaUGMS8dc3x5gSjCMxFijGOr2y4nm+ZL3Zw9wtagYujY06IHFmagplwGq2Z+1ZzdpcE+WZ
YsysddpPrOsYGVIdoAdzkoCaHMGdCvhhotwJ7E7sc4wDAbW53P4gkNcV945/0e+z+NL5l9Nqig36
xU9ugHoQnJkeUZT38tORRI0Y8+odbUCwsOl/54JF+J2M2N8C9HoNR3wbR4kQqfWrPdvZG88ednDn
aCLL4IIZmqVIdxtHieCTF0gnjXsL698mwxAGGwsbqPICsBlCXp1gJr0v+v+dzYxz49NSutLDFiv9
cPyuKnKc5iq1ey1c0GE+XMO0n6XttlbiZSwRJwiySx8/fQKSxXWKDDfqCL+GpiZk+NkVIIhcCPGg
qaB1pv5VlOxG4y4tE7rcNOwC70PG8k+ZidavOkKyaBi3xq2rfmlilyd9IvwOCYkuJ2KH/4uiE2YK
NTAe1n3YKCqcEDEbS8n0GJkOCgHC2uolRP0i+ENqD4GVRJXqQqt7p11rhqqcuUDXTB7dDbPER/vi
xkrSffF8hCGCRriCAmCektrRAc3iK7ZZBJ7leqzK4rHmcHDzgQ3tAtJ96fFN+e2WYN2AxYNsUHkM
Tbzy756pvClEnpex63pFvU6eBQt1nRMDFmwONbAX3k0x+DTXD/VSgW75WPKcsuj1yX3uDlvonkGW
39tDnj/yyo+ECAHqeMdcNJIT7czATrzV96O9o6JXUwXvkLF1MbzJd8gmEb2q1u5SZXg8reeY3QoO
t8qmqRNjnLtwy06D8ycXrSh6SU8ae4c5IMPyaKo6EvXKbThjkrBtK9DFcinBFeuJouTp0Scxwo0g
zOmF88TBccYd23D/Z8KfCoogzFs3FdyDzXkueSQFWl98UQCDuP2NsluctWcxcBpH3QdQB6emiZ/m
vVpTabOW5R3ozgbBltifLbTksNJ4thpI5ihzhJBS+ZbCgRfT9FLUn4Be9ehy1eIXuL8cZ1nzWsGN
gwVzBGF5cfBlZVNGikHZInxYmSFvENRTyAyCa90JX17l6/vGfWoaMuJQSn0HY7/NbM9gdjEx5U92
ctDl8oSenTAb6q8QESYGMjOabAF9Wrx6EDT/k0HbYlCnt+sf4twhzqCDQNXr3dqKoSxm30tOUh/B
vaML9sqlcYEpw79/GZxbxUuU8PdNRBMzoK5RPoBS4xLkJ3pvvnnqFzCLSW8biFtefvnIIip0BPho
eDIaACTlmhixBpK68ew360wswAiG8cSFX/iPsYZJ2XTl2dV9r4imeW87I+T2syhclIkFhpmceRZY
LpfuwV/jD2Hso/1q0QZgphos91ovdxh49FgujmrAfkyhWv2bdb6JohjHEMmZo2ctzq3EbpduT3kT
JNk23MKOVnpbBtItaRhA7+IguFSNC2kkunIJFWbdaItqlBNcIu5894uFvuIUp44QQ2qVoUvTMlcV
KCYxiqn0elQwNO2jemo58SrSOu/xqX3tc3z7y1VmGlDYPlDoSYYIb301RnaV9VNSGqlucWyMlLdr
VVWDqQ1yk9X6iZc6tCdhGbk3S7idWvWiz2Vc/Ko6/vL09oYSgVcTZd8GU7eFj+yGM3q4MYxUZf0/
04TsnfZMNw/6ZCQgI5aLZ7X9D0dfaGPoPNS22bkosytlLlLvYgi1gzxjNrIA+KkBcqanlWDPIT2d
ueWlx2y0ocYK2lSXJSjjiaZ0AqeJ3EB9JIHW8e+gAgT/Y23izhP50IAlXvi34VwU8nJ7pNfAin/M
NOzZlkU+vF37Z4r8+SO2x7ASfF2OTK9P3/QatbtNkIv/fBWs1FcDxByuSkV7pr5rrA+HvNicQA++
cCRdn9ynnHK2UCTDPmHdgEoN980RvJzl+NRWBy/GiG/7uzFVVmgDeiX4shKyyUp+HmpEAv8+q8S9
/cu9d78uwi7LmTzc4wp6FZDZFy5lUaDdWwG3tfCjpGuI1jSvr/lu825B+ea+IRAJVmxIzatqaoi4
y5VA4e2WhQF1Dn6Z5/f6yy8SO4iCmkGmOfEZ0yJUMtR2OYhIjIeFTpLKlyrhvT/oEsrJBSowciFQ
UywZh1762fRJKG8pw6olZNUFrKPTeJyutQ7BKNT2TFYc1zSZqykznOnpW5WbQF4ajXdK/z7Hj5Ox
Oq0YmREJ96cQonKU0iYzdW2qhtH30YC3d7jjfXSEfNzi/6YM3CiJRsuvHwAV+j2Ve0rysPl1g7BF
Xcn0devoctDf6IGZt5KXFiKXRIzLQDXQVB4SMB8TDzGqNdlFRhiUhvC0ZEnjsSnps7Mh1tH6eiab
W1v5QHs1VBeIpQhoAftdwO+YgkVJFLcsTOT+6oTX8cxFgEn9/yq7mH8GX6LipMWD8CfiyOq6D50b
uqCRYxyBUlzFHD5aRU+8Fv11c/qHkD7GKkuSepW8Enq6IY1JuJvHkCKiBngCUSNBShVJNPVnPqbX
hiUEd+8rdKcA1iw2Pc8mQC5XwRH8hHGeqW7BEkFnKTxHlE0aer7mP+pkFL0/ErSFQt8o0SvIS6ms
bMRO1IJsAogiKyVqvOu/XTk1oRyhF6uCJ3CFlYyMvSIqEAfk9yMjOdCi6/Wp39JLAm5iZAB8A73P
Ci7/ARgIpuheWYNYyHZ8PwXIQrlJ++v4UNHVAUbeCCNDSeBGQDql9jx2uCZ0nMpDreGILVVZvrud
8KO+dFbtR2fhAunoNSqisQOLVeBMIdVo3tD/i1jBanyfk89uRq1rz9xh5bCA1crr0KuYMvVRd0P2
X7oYtRXNVNYCvXIqPfr6ZttjIquQhUxqMbqnLEHjlS7m5N7yrnu0VMmt1cUKHRliLupS9aS5vlmf
jgCA9MzmoH0hTVvovgOm35hDlrEMWZVyzrapJCMIEVPeWUf0alLlITk5h4cTX6gojtKs9h16sww4
fa0S9PDmNE1PWYOlGH6YOsmCQ1Lj02efB+8Rg1Ji11mkFxiCbvZgsQ1BsmncIL/0Q/fR7TbDpQIR
bRGsBkqgTvg/Ccgw2DNqyHtJR8Y8cUPCFjWZ9vhdIfStZnVYuh/UcjSGrDvq6tiSQEhTpzXrEvPB
nWMRKn751yAppQ3qIrwYTLQbDE4qY+MCRM/q1mFt3DWvE3r1wyUk2d9EZz86l6v7EEIKkumaWVn+
yjj0F9ES9P+E9MDu8Lr3cI+6nOMfwJv5kqaTg2ALplQj8MNQH8BuVXFqk4jwyako3gC4pfspclMT
EfhmvA9+lgkIVzYYWyVPyG8NxtKKowLsjVhtLJOiPMfIa/xAkT8uLbpQ5RzbAIuBfdMskjZQF5P1
9qKToVR/XKxwB4YV38DPguTJaMU6ALs2WQ8URpZcOq7AbU6IonN6LkRv0EHuMU78mZbMM85SP5yy
Lz2jtfcpgTZ0XDVK2+U9rlv7HsdtavrMW0IrXxOqUJMkcx7s47oroT2hLWVrSVGYBdzB5YdfhDRD
SCEqaz/C/u0up6qeG+nqfgTB4d6Hgimgw/a2jADY4WneiGR51dGmAIOY9xrvT+MkrH1U8t5eP9Lb
0a5k2Op8D2jKQQd222bfo/DZ/0IZoCDHdc1fp+r1VeeBsc/d8Ez0wiTPusFefAGI0mZVVQxQIhza
ygaSGQbOjjWgKCpsW0iYHTAIWSpB7pR2TZdejV6i/viBSyHywJkAWOLKe5Mdc2Y/PJV7Yg5sBKJT
hM9+oPQ8nLzs9iqi47IeI6PfjDTDyt1ROFuuWVJu1oifonUs1Sh+KoidpipSA1m84bJd4Vvt2ZQN
uZa0SIjIZ0Foo//lfinTCr4DNPEIOee+ZEl+AhWkvrQDiw8/APhA6EYDlKuF96yk7VvT4Lq+Tc2C
3DlTg6TdRE/D7cFdUYWDK6v1nz3syPCTHNYClQ0GS23jagqxFDk8n+nqV5ASazEl6nw3CDoC6xIW
dnQDBBlP7eZkXnQGCd0spmIO5+7dnjn3ho4na7D7MPclpGiNNu6PLkXwPlIpAbjv1IGglLzplW56
boVdXNYGXwgVSYQbr2W80m41xt+ES0ML/SSlDI0jgZuhvzfLwdCZx+/Udo7haszbPArmvwiu1VWC
6l1zq43hHh7AOINftf1dwYTrlcurrOkkSu46GdTKNkMbophyFBP1Pz0jnzAB4jckJpDf9UuCKq+V
GWTt7rdb4jRy2jZZmMXGuALLTdVZ0t4aZOXMiwmp4bqHVX1RWURyKPPQ363ICOJqslA/1UorGBY0
8q2ycCBgxst49WkBicOwSF3ouwqQCWyOMv+5LDPWEfcEotwjwNdx7wRVlqL5B1vM28FITMv4WnWS
pHVnvz191AguFk4fqt4oqx+8k0TXVHnkKvVw4iEcU+JbQfY55kwIdzJhjrPGG8xPJuB8WUGaNSDH
x7bjj6lOy7lcd/cColTDXBTJlS/pSpq1PtJxNH+wdyHQ7TAfFcoB8TMIn0IhVXfOJYZYLqWysIZQ
h7giJ3QWKgFUDz3QUqrqByvT2vuth0otVg78MwN8DG04oMti654ON1ahzrk96ykfc3BGbWFBeCso
twfxdkbfUirHSGyv8ZDEO/ZdozpkzL0KJnIjqAZJoRFj7s2YGSietJrwVNFdEr/7rih47aegTiJ5
lRMQc1QVv+09bkT40cs8jHp2NcPzfwxldTKZ6gdAx/PZ/i2aumMYHVLOOe2Lq9KUKDDPZQ0BDrqt
fDslqMV5NSsfNYvuNEpWwnzbFj5DuvEJx7v0dcx8w5Tlu9f3GW+9f3sHGuMaUC4c+b74BEV7kPYr
mRRIkiD0OUMqka3Wvj8vL9B56jeRNEmUwy6Csv5u7DXsBA9g1G2jNuPcQpTpBtBjinS0ynkDJ6da
LQtwWqCWTEIuOGaF83iqOp1ASyGrdR/MWnxzHdJywldevBeZNvx0JvUDWLlKSqwqbtVhY2ozKv1y
nnBr+WB0uWO3Yl8iMW6wqfgQd8C4Nky2oHAiPe2wDmQDk26swx/rYfNj6T6e151zMqm3X9DNjXSl
i1YxVz8llxx5GWhuRl7yu9TjGQGCf6uqX0nwinTbwo28+9kREIgcMuxhzujiKooCjrZYSCA9drgz
nKzrfU89+U6h4bo3dBg4c6OGQBnzqW9FWw/1AQdBOIfLno9ruQSAI4SCQy6BB+dsOTD3q6vlraNX
O+eaQq0hpkxuTm6ujoPGXyDSXULoVaLQ1CkCffiRfFK5HvmCk7l/StCRhpfeHJD0S1+2DsBkh6uf
gQ7hroC7IkdvaDtl9u6SB78gfJUxE5fNgvOdHzoqiqLPIGXi2ECvUfsp0ZOJhmcBI4deXSKEOh1a
+lmrKZ3L+icNMa7REqy+SqEwuQRwQZqD1VHYo6DBmG6uEcT9FWyNktFGrv2lIJK2qL0i6z1wPQrg
X4yaI0kmw1hTLdbVTaRn//HezFO7Hz81IFvBDA2dRadDqPoo3WRMCPh9RkAeFD7/A8RFOhqp6VL9
L0+Vv0aw/J174mthc+xM9W9jZCQjfNZxQigCBy4rKIjYxtOETpnfpYkx2Qx9WuPaGx5itYykzL+R
ebSzvMhv1HQLV9E+TNbjrNj91oxFVkykpKZj++jhPPHlTfWefmBvW3hZ2pvwI/RoDOsMMKnggfre
0R3Qwdtzxl44pL2+LLc7jJExFSKtF7imkSSVrwtezq6AkW+k6rMS4UU1aZJ96S2BNWllAKoUWsnd
dAOGCi9ADHBg2HbEZ0Ts7xIeo0FincQbSHte3BaA9OrckCjU8j2X/gowBQRs106J7PY0YJtWVCpN
jvonM72L2bM9Z/EUOUlYnJOaT3yAuMyt50+fRB9Wm1dftHW/mqtBJG0L+1bsC5VgLM8eteU3mL2c
ofHsIqYNfyYpauuHhQC/b2va+Bzo3xSthIsMAM8N/69hQzX3dkJErkvcSm/EM7YgzXPWvxxFNx4V
o2lGdQS+oIpQkqTZ4KwarUhbbdN2REymSKQweNMpF31yHGXL6ALNSrNPwtaLKzsxoZrSmn4If7Sc
2Eg3iyTZsZaKOxQ1gZvOTnS9JxlVxT+Gw0uK4WD8ou5tjTwzHxGiedjNv5WcWr4oFknLyFbBpbwV
zCOqoqkSc53sKGRkRThHvK76+HbUoAH4Py+PXA15Zg/3SMDEBrQqI6a6PzNb1qpWHLPg0QNQB6sv
8ZI1W8+Ujo6hhiVCwJbXsdeAp5detfImm/ahS0lIQdS7oMnX0w+FPfs0GHqXjNIVpv1mnxUjqdZm
gy6B4v7QuVidedVnGWjRh/8TJtlEmqAjrIBwTw5ixDP7Ie3K9dH+qk9wp5YWvn4AOtEnNFzQIMac
EpAD9SjNzSDTxvyeWsxDkExFapCFmraoDUwa16czFRUPZqLDRmYLcMGz8CPfrVWwtmYnMrwN8UiV
WRjJ7I77lUUkhteR4FVvTD4XeIkU2RJilpKwpu8Q6aRw/y6Kg8tKhEwrlvS0sC3rUirlsIc3KMbG
sdIy4rI9ZL4T4HUeon0aZo3C+3CuGgF6Xwgt8w8tw4HnUPkobsNAxzlv471XO3nWOXB+ANzw16M1
JM9QPz9dCuj0vJ6w32UmvvJl2hDubPXtd1h0/Ro4+kePkZZn3Hv3LEkVXag2cOMzVK0bkYtgPi9h
BEJUk8mPAI20EHZPuVydIHGHj0eCU8ponQxVGHfUxec7wuwW1buDff0vyYTtVpLjnG90DCuX4xyM
biCkGPR1mSWbrZTvrO47qnR36jOg61VZlaf877pwqrCbxi0F89vntCkJ/6C/wCT5gYkejZJTsJbw
M/lLn4C2041zeUYcOmoGcKr+mJnhkRKg8qNNHoiDePfP004QIMi+gwLS/IhT3PYezXaOUNAwz1LU
ZglQvsInnhVhrYdY5ogJIcUtmmqkDgPdONlChDXH6LcI1Rwi3JjyRTH40rNl4QTyjUCu3A0AIUlK
GPj/qg7p66INjwlxmF+Z92TiXMKc+cwDFAXK+NZ1BZh04nWyor2HYoNrLzixIoUNWwESa4tnSJfd
v/ZkK13t+/K0c6SnggrP5q4cHdZVjuE6FOO88P7nbM9Yw6ubE9dS50Jjoja+YKXKw6NltNB4tL6w
fLYyW3RmyhyII6kYtxAB49NBY6cvLx4z/chypX3XnjqRg4umq4Y4iaKB5R5jwUqRCKwo+P8qORqF
AKAogYkFfRIqjcx3PKRYjiIxwbSb05EERDwVLKELyZeU4nxQUECgX+2KytpUES0YFoWBhYt+8/u9
J6XpUGpMuINmHnQIEbG1NKmi7EKmEwy8oZZJdi4c3ctNUBmo7f+a8AL/DyQHBQ0q3y5YJ32XtMz4
YQQbadJOKr1OAIzDTq1plaPGS+j9D/wW2rrlQjf3Db+9ILN3JabIIHE6jIZ/DWYcS3CfgvIsSQmv
fSErcY+TojSwGifGfZbvsIYEYoxnaLy7xrPGuZ8phVCoflLdbD1xGNSutwy/1VpcwVmkNHGTFinN
UdtN/RJC9LG4CLuBEjCdnw0aJhrTQ5RoJ64wQcJN/8UCmhU6HEgLZWYExH2VzrAVQDmQ6IRtWOxu
DobB8aHs4dcroTrvfAq9tUjGuXj8um52AhtZMFiv7vyM3/RkPDqj9G3iKeEI13Y12ZJF8F+buKEu
Dv0yfi44cI8x3J0z5l5BGkaekwCvvigA2peAKo62RNaynq8axmo0aPS+6HlDcqXHSqImgJypz3dQ
n/xXch2Q06XpaYpOd6hlll1l2f2K7odh49qXy84Ff/5EIpRboofsW5vxIfyMXlMdwVc58EEln3rU
7TnkUH2C70Al77Y44AO8Hq+fWF3CkP8/r1cwIbdKmVYB6Om/v2qDkfrdF6IctATJBjusCgmE9kEB
4eSL6gulcDZNdJXdRnuL9L6EFawys4YTKxSn3secNCfW7rsZclRr07acEg75mJDwdk9pkxc6GFEN
RWuxSs3usEVAOdD0KwH4LQg/nz8/PGkk0q+eya18PR6aJqMgtqEZvKwYPUj20Y5mu9nUrNherusr
b1/L39Fxpf0tX+71/sAsGZZsH6aP0pyagHUzlK9mEyxOBEokak/h20l5/tBaV3ZYO134LdDTTD4Q
0KXEiHW85yVeCX8llSYrAKZBTKXKj6jQAFcGdXMhiUeBmE0aJY4TeeiGVpWP8R2eVNFC0S3u1fkB
L/cZG+Ih+23tB6gob3czvckx9I9BOne7WHFWijgszd6knPRQMKezDwd6OHNlXRnFp0uQG6C4/br5
D5BvGIbeHtTAstGa04AXtfnl5B/2O1v4T++TZumVtFRqdbMsGJrvL/ops2Kke9JdW9SRJCOLF5v3
AD9ntW4oCVyxk0BGRpFab46oLkJstCC18iEPBw8A/JID3a+E/MMZ9N3JnJd6xExVq++U2XQt1OW8
jFkxPlFEqR+zZk9qU8KHp8CUeVCUIglit7zsHDsFVG5GFN+MRHpCrnKLYRuFmtDCjnVy6gxFwJJe
Iasg52oVV7HGqaKJgjrcv0CVVadjiQp41521rKXoieS6TlFGTyATKThsTya4U9G9uc9f5U3tdR8X
yDwaLg+XkYBSR64yFd6Mf6WIUgWTrgit/0xF3iCJYw+d6BkNwtDQ6Mfpf8qsnlbDzYrgzd8qal6v
3BAwnwAUMYBE/tYpRp+STU7UaV+4YHhhAFXQcgtQnghmA+0uCjGf2Hy5Q3ZrxNltu2WsbZ80MzOf
cz7G2Eu3/gCJX8TcAlj8uerlBOUdyAWL+Nk6Qn7ZQkBmJJD9yqPuPQQkhrPsLhcWWRKJjiU9+vVg
DD19p+gEPQsEEUXMyIX2RC3HIyQIfHPzVwUudD5uFAkcP8F2j/LjvfpjW/EXNQRgkFSPpcAKFuLm
zuEWBKwcHdB/0n0QKrfUjnBgh1Apj3Ij9BYu5ImNKLKVXtkZ5jgLK1WgDfvKCasT8H7BBpFRa5H5
Z5ZGORE9fEm5PK/fCmob31i71KmjsWNh7giQINXFSs39Zj/OwC8dwABmCQThLnzjjvChAKxgKtSN
KygfYqTCW/oaNNSHRqbE8qWOYuhpPlq7QmOX5/kOTJ4fd0T4pSiXnw8Y4gY7ZJiMa535G/JOFCgF
WDMAoVW+HjHqb+f7Kdj0S4P53skBrzx+kW0BIhMP0SU1hpJeTlMTDoSkqE6CQj0eafppWjfk186M
cjaT6TTsURx0RYrf8/BW25gFRJ5QTEVxtcVsXwdAq8j6ooHhP9FY85UL1jS6gNBbuF6z512nJ0cD
KBpGt/BPEJfzCkg4I7hSur08hDjvDD1OFw8DOWIUiBSrHxR2h/CGW557EyCnK2uDGta7RhjbFJZk
/STQy8GvqKZspxj5NWyCvKWPigvm9YdFtsuj9+YIxHGRfKWgtYnXyp0n6bZj7v5CqBn5pRBootBL
DypnAcWwKOEadVjEMjj8qE1TdiDUzGq+Iqv7yH9/M2ScXD1sstJJHCmOHzh6MNd0boKXdd2syBQ7
rksIXlTsT4am1z20jXgcZgZKhNo1s//YRikvhbEtfq1wkgwBvMrbt8vBmjabQXrQtWs7XsJl/iLq
P5FWsS5W9J3xfMd5Q+4EZccqa8sI7TwWNodKcocGfNdGgwhY60XSBIoFy6153lCZs6lYqUxuzEwK
EI3VnPWSN+aBD6wKmu145MWOn7+I3HzwOrE1l7WYOoBqndVPrV7XxLu+W27PYOSejb29DdBCQ/kt
yncdZvPWlFF9Msn9HHzOwpQ5z8V3e2LKokEl/pG7PuwyX/VLunbEGn9NUlPoS2DLEasSHG1nUOF1
x6ZCrEw7shawptn8FU4eNi4flk+ndFxoB0wGlCpzTrsy9K64DUhkCqkwEfrmjDSH6S2PwDDu1xsh
4vr5N7kaYKxi0MBHcGBh8C4dk3k0PBi+tsF6bvzMdCIbOfnvZ8oK18tBvBWCRe6EhOEuT/h3ifbW
M6Pq8qhR5ptd1TUYOWhdK8rza0IbIt8Wf5mPA/9eGKV0dn813Audg/iVosTOvXRHVyg+x0N4cfkh
LV4yK1u++z3VM7yTVn69ShZ8UVJLQtNZvNSb/P8GvZAQNdJUPmqHLih984le26E0y7A36LuXZi7A
QZhfeRl+3FOO6GrXDHkuFCLJRoG5b+ybprHXT+CycXdUiOFvKTyWTAhEBlt/NVOKNUCwChL9j95n
kAlCMu1czQiXH1ZuR4q+LoR6xSika3UQScrlUrVsLDkpqGM0JIDewwcq8gvTCI9qr+tjxU0OcYac
tAfL0EUHH9h8ddKj8dgzvslnrSZCKfTwo3NhGmqe5G+ATMkE1OXcdfuZWYn7xH4njuF2sycwWDxe
Qq2VZC+wSswZU840S2uO0nQ+kXUe0VL0zYf4fSYkc5DwFwQiAnIOERfeuBVCKmgtu7dW6gKJhkZh
C9btcnDPiOMRyrMcPprE0HcwJUtY6GMRg0fpSC9oYqon3iN8eLrpSUhfGndt3JxEYjuIxA+cC+bL
7HV6eIakDq7v25yP1H1HUZNOtdo+T24jzpffHC3SHm0rbus+xbHuMRe7hXgJMdGRQtqXAZ/vDBxA
56MNit7b1ec7N7aU48tCs5aHYq2AHlxxTqcwvJ6xfJH7baIzJs/PzYl5gDe40nzwLO+4LBt6dskH
hvx/tmqR/lleUtKgaOElAmq9jyLTJNRBtmPWY5s0Gat/xIFBaLmmRpy9AJqGnQSJDvmzdB9NiswA
1tl2Rdc5jNkCk3lM0qjOB1TDpBFiVuifqSoSLLefBW2npLaKa9ansc+m50wntiSwsYb4g/PXac4K
LJ/wcVi3JUB1DecQ/2p3zOx5zl4zvdkP+4kEHKdIg94xHfZxF9t2CB6FFC7Lc6jqsCxX14uX/Qjx
UT4PcjUyJPkL8QJxLBars7Qzj95DYh+2FPa07tfqtSSXiVaNcGzVqGPuxsJHP5FvLbGXWcGkPgs6
JpTc4yX/SpKo7i/q49TdxWjpC/1Hnp2Q7uHxzWUh/U/+0aZrq4/pDmXTMEeu5CyMPaKnv4LE61aC
zty4EBpJgpFlbs0bOMu7jKBxrz1gnLUtw27XMC3YLHs7SAvPEJ0QnSrtXNMUR7fAOB4dm+cBeQ4b
xVgkCF8vSZw5cOkaimNgLiqOBpjc56Dibsn2HvHBZUhBq7ZI9zSsmhGpVTq7yq+xt25TCwuLYV1n
e3VILv8CygQnwjsMjHWr11emGu1XE0sysh38uabb4A/GKD5JPnUrpHEe94JmpsQ5MH5iB39Mns93
svnMAFnlmVzf2Mv66yVVJowp+xrLd33yg4b/BeMvzfAZd0LBzPFDh+aUOpIER2mLmi7dGt78YzM1
KYPGfAgwYe/s1uSG7Bq5RiBn06uEgRQgj5e4dGrulVTElja6tDnfxD0cuTbxDUWVDL/03z2O/Jg0
/gsqJjiW86fkbSJYFLN97L3Yd6xOQD6iwhIg4iELJhvzgVGfp/axIp95qQzEJuuoOUGp1mPDP0BA
BjHQNoFHUEPIxxC8nAK0OHTxZFnSs9MD/bCIRHdIgiDOTQsElsL0fHTckS+C36+DeERF+0cBxGji
0w3LDCSNzeuUhdSxg6yf9A7Oigbk7GfpOp0NBFib9gUVmuvng53AeS/WxXiGWjJmmf7MCSTwDMkO
8Ia3Gl8qyLWNJirnpbegJ7zawkOivVCmiwLZT8lqDvzUzuX4PKSsqpQq7IfFbbmXFCOiBdwt1ZHI
4r/whoVmGLipFYw4OkfUoIpAyyWkOkSmO0V/LHqzmJnZRAbZqv9w9FjGSbCAQfasLQ8dJhQVfv/o
O7huOJjH2ss0ZX3IeMqJeLyulR9Pfoa9HURFax2RSTma+jCNFB8aj5oSGHmficdL1NFlVowmmeKa
sqOkUi0Wnvg//5e4kiRpfJn4Z2oXKMi4RHFoDhpYs+oV/DweikIVIPjjmP7PXRtpSG/zefrJue48
78seKqiPbRlZWgSLyXycC9VZ6DZhAx/uQDTUpmJ9Sxudw+sFLO5YRO29zi4IggO5D6I/RJshlXE4
siF1tRNNf8m1xA6JojvyOW5uLZPLYrO6xJB3EFDRzyKqqj0Y5uUvKn3mR4GpUBAIyVNatUBOxNhc
Wer7O1KYTpBsCAdqU7TvbHftTvp+b4b73qxYFjCxsBCcjrs6N8jpLezEUSzLX3pz7A183PKoLVsY
5jUoArFCBpJZB+036OKkw3M0oJjLkaY5cvDupvRy4+en2mfyTsOepPszRTMkw3U8hyM0eQuqDXWN
xXkerm+bCHWABngw1UKi9KptM5EW0S/CQByb46g5ee0KtGI31IvR6sIvQdtapWcnvkvNow+Z7wYX
Vl/MZnQqj37wxRhAbhdM9Qa/hVZkl07GalEedAuGqWA4D8/Io2EZtL1fwAA2bWCv8XRsKgnZ2JUx
XIOwIV8pfV1EXEDk5/8N+rcXnmu9nz8wqmY3MwEzm8cW9AN9ZscLrrSa/HlbR4fwxVUhykVbjvL6
44KmCLlA3lGaccq7t1ARaEgXB61BQhygW95V8RxcYV6egCqKxNvqCcQMxOqUV9zc7HA9eueEUcJI
oAUh6wGDTTvgZ3luMQYKBIgjPE7vEC7CAwzH0rs4qVzXszXaLBBIAUsxqERGjxOptViGk2gl1npC
H+4KbR/6G2tFPDQfUnLQXfiY2J59rDRb1iLQOtIwXmJkgrqJ3OeAGZTqpTp7c79yYiuu+TEkUB2i
BhYKxdpzlrl3G0XUWu/FSI62dXGaBplF/nukT+fckKlx1a4vgvCxQ/LrBKkEH9DZJR2MXmQJElxP
p2AGZu/RW7nKI8zt0peu0+DuIQT2zdZ0JCxHmnZd8v/cC6xtKytgx/Wl+QaySBxE0zz/cDfsIPou
h3JRtoV/A6GsjjCD3On1g4Zo6iCr/Bw/O+P9d0uBGk2Mpb4W7JJmTzuXfb2H6+p2OaUXU6hue9Ch
oYZ9H/BwqtEEPJNwWXnkZ9qY2XhvXyJt+eIFeXT5TJDJzi+NxgUGzAzOyK6qrrq2C6j9HgUkK3J9
e9EwA92kHifZkEf5VmgEH/Di2V0luCpSCIA5I1vSoIutbWeM9UQtgiHExdO/GtrNdeT2cH2dJpAZ
Phe1JZ2ABfoxXvnEclmc05VaVLHseXXKq9oKkfvoKMwo/roRx3i6yHAUD7tFbtSOqlaM7GmlG/T3
dEP0tAhGG6iUKOF9D+qMUJiq3dy5Yu9tzJ/HNnecQvk4H4ChZ5Mcika1jVa9ec9j+FHtJGA6B6Y0
QvI+BhKHnWL3InaJwDJvUUerTvxG4JasH6G77ZdhT4H/GoOjBcEOY7OyauXJ5aK25LhYDHEAHgs6
bM/l2u+5xAsn7WQapwi7DE2NDsfSD+aIrEBHNFIfrCQDEbdPyA74NQMSQyVTCtNKTx0phzJzEFHc
pHNbPDvrFP39m+wqsl2L18dZ3mikmrI4aTp+GsEpTfRQoR5ZMD8Z0TGUK0q8yZQfS780WANfty5M
oenEhtEBn3JdsARBHpxzSuvd9eyJlX5y5yw4V4U2t1Vi63Kt21NgoTuqRjS8ZCfiol7QSPoQWxSI
1GH5K75ByqvfOozJV11nnww+0SEdriK6NwcHvhglqw3GtYvx3RZEdMyluNuPCEwRYKoTiZiJfcZa
sT3VeHbLyi2GVnx/WbAPzPvmaEd40yQg5+T6l/IEQbQ6hA2OtjoscOhk43DDNAZ8bFgx5OJONwVN
RqwqGo7YRbjdM0a814ARQ5TPDCZr7D2UN/1H60Oh6GZgtO6d74SVHjznxaLsGsfnds8JqptbjVp7
2ZgXd+M4SM10nweCI2if35Jl35B8Q4r7ERzrYWXLNV/e3J4bpQrmIviwK8nVbcw9/sBZsZOBAdGV
7LDJTUtu8r0iEuvpuD9MYpFCCrTxCOVssUtsH7loo90vHNMgnGJ+/gL4qwKlJ8UPoWfcMQWj4eL0
Ip6SsH9zD1WoXwu0UBhsjf1QLN0RXn3pjlpyZcVj3TEAJZ+gwG8iXg9IYMz7VtGm2etZDhpE7D7L
AUiY2Eynh50gWjLaU0nLXnwmgEwsa9Y2Void0ndugJVy7RiV66yokwOaZkEYfgV2xQCCZ1OIphKo
X4PVtQlQfu7LUVXME6z6UnZOGo/lqQuteWues0yHVNfGMQpe3s0cYkEa/thKvmjLS/0f5GrQ8iAP
+yA5Po1QbnzSL/TCmThTXtQmunnovptqzcqxTCFhoiQvC+9a6HURIBSZFO8LMoGoGGcjKiN4c96Y
s92ch2gi2VxToWkPugx/EyjQv04OLGVpVa+WDj3A/Kb3hGTseMPfW6gc8pAWjxlwQti+K2sBEE82
iaru2Q3XipHXOU6WXXjv9gNv0Eo/L7DIMHmjfs+/DGIC0SCv35tSL5bkwolLEcNV4RiY8NhLYuvE
JGQA2bVDLQryJzxwIb7nMX1H90KFR8ygC0zkvMNZ7jD3a4CfMS2Q6JWPnVoMzBA6kfzx7mThHQ6P
ajRNwGnlFQB6hhw8T0dpo0xzVtEMAPBDq5EJCoRqhSeNXMMpxbQCppraVvVVu4+luwOTIn/2iOj9
CyMss08XmO+Aiu/f8oemV0nRF/PRcDhU6MuNOB5pgSROOnF3DgBeCF7EgOeTV3weMlBscOAsfCZk
qJA+efFbn3cI1dOHKvAtMOpWwRjybVn2fOj7gsHrkxNDsWOFDkUYXw5H29kPKK0+H1K6CSEGLjxK
hP2ZodAIrlFLBDNB/MCjmE4p4LRrlfk5BzF24yhECXmf1QhVcqC3eUyS55rPAnteX0WB2bHdTtGm
gCw835ATamp/sXLqc6xrA7afOG+pzAf9K+jeh9oEd9kqwRAvuk/Mb8c9Jc125j3OVNU/na9bpJOx
4923i+DWxZYEX9Ta8IRD3vevyF3j2zk1y/Wqe3xY/QfIMkUT42raXbbW7v/6OjXu/DXlN8Kt9gs2
tKvqpbE1hgw1UqOjfIpmoDOASkrl+kOz9nb+6Z0s3FRks+/ugf33LHCrklPp0zICmE1OT2wkL0BI
uNXvwKvZ5vAQeLEAbWJ1KQFdV7XAIKDU9btUyuwc3r1DiIE8mcBsfjFTm18rTHGC90B4eFFO3vIh
dXU7tYdu5FqMu97biieKN3bzDvhneG0AyWIbC3/4vQdT52CffDulnwag1xLCMs7TBhHwWS7SYEic
/AayEKCvCIrPYSMgk2PG1ZiAG66676Heg7GZbtQjLQd61z85dcQuhKZ241ft1BN0v8/3Xfak6ElG
emh431BCrJ5Z4EL0qz0dK0E8PAvoobjXve+NJMAtAmGmM6FV5UybZWMOJAxorKBtJLBmQKk/F0ya
zcI+sFP1XGKOOm1BuMZAIaJ1yILhG+O6SvGLC9Cl5lp2rqGhKu5hHRokf8R7YXxdap5WncdX5Xrd
2oaSc4qSB7ei/fyvb4k+Ba+jGsVmyEZXCuPCBfTzpTDmguxYZmXWRfmTV5+ONmyjj2obMnqMZ795
n3GoudXX6kZYMHmK4jWqKRthKleOPuGMCe+2K/rMwjQRJprSSlPilk6q98/t13cUVJLiKIo3j9ZV
Sd8ZYtEUiZzlanvqHbvd0chXxWKnOEPuQOo1kp7Cnwsh9YhRFeA3sHgupUe4/jKXo+Ugztmbyv5U
/EI4iXX9ubTQDxJz5qAG/HNFCJh90T3WJ/XWUrf/2TtwYH+ijCbPmYQYej/bHX0rnlS7WFfdJQyn
tdu16Olq2zUlHVcyQLf1439nlsKBEM1uHPKH9iJhI4mO2bbchzbrmV+5IFi7wL3zWvq9tfa3zOQV
muGwWy32wEhtfiPiXvCqZRdtQ30e+rty0S7h3aydFlKpjZE/mlsu4cFj+nZOJvauDIZRMy9AR7ra
6C9Lf1j1zbzPij85olSNF4jifnJY0VdnZPrAe6iOop3d08rWnMtqA5avhIbKNGlaVyX/P153arYP
8HFRyDKtI85zuvMf2ALhaLmrDQFphDYfWIvuDrM7VLmFqbSqLInHhDQ08fJxdBUAiYDeuhWxqhD7
7Vu1fSge05uKffZ4vlILOo+7dMw/BJgoSvddAT2C6op+7jMdwnDjGQHbr/KeVdnVa+Cw37Xdgwtg
NQStnJ7Z28yc+m4NSD+GB5WkAGy+ekRkIcYHjl925YEZmDq5OB2LNaZr6Ffn0X2gns+FL9OuJK7s
rhzQ8Xw915kwAHupf6OCReGI5BzfIFthBx6qtzCUqOiIc/U2l581+Ss5oo0JZIiar7demG3yvx6k
j23OKOCg18KqIlY/FUh+0AjEVXY+dSxvKQel42wNjtIxTL8V4PFHKeroQe7/18IPg/zGhETukEM5
4AtIf089aUprsF5k1lTxXaAiqlE3oNMKZn556AH62ZASbdF0fpLVFMN9SzOJLBza0JBibmxpKosu
mjzR+noLwhakUiAdF1LHCmZsMAgpQY38iuDv2yGt3CX0SajJqy74S7LRBV34elvNdtD9DNijMs5M
eBUtO1LMZ25BJTQEwKczrQV4t1kz49/zFZkP+chJ1omJ3n3mlxxpYTx/yg7PWa4HudVg0LIOf11y
ogABzLCl5RfmTp3K+HcwbaLWVB9Tmrz1+aKZDAnZ6E+b9HT7MhcruisBB80GD67tRM/eSc0ZVMZQ
sLtb/+u0irthpYkwU99eUlu1r4h5wnsFxMCuXHWusCMyPWBavugfOfxDJkuksd290Ga4VXShecRg
1BeS2A2CYQ1r0E/D4oiEtkC/U1arAonRd1rrsP+KmVM9zbH0DJl6QEmPOXt7mII3rT/0VlrxtKz6
bbrinPffk+tyoSOBkJjZOlvFLK3BtNae3Gc3/SYrsKCOsS4Exp6CAE20s+x2PkvUCVpuAYzqvXLk
o7gt/SiLv82kaCRhcO4K0CrIbNGAjNdmSf5fVu6FFEzd4OKkgquv9VOa+OAQ1wTIXtns+Rr3SGQ3
tdDuTQvrFqCEGobFsiVJ6ARjax3dv6ErYE52GAfWkDh9VYGpdt/+6tLMph8zDcgRmpKB9lXZl7Yg
kLiYECAMI/lGZjh4wK4uAIecSTr8MkW3oM6AY0kMNXgdwnGf/qi56bd8+ZKzlsgq1951I9cmQQhv
HN5MTG9ayE8rhKHLpSG534WTzqwN0pKTqfFaDZB6Dnigmfdb1JLTOeCCcTn1Z+UL0c4Y+C5ps+5T
G3JxWLwZ37THe/zKol4jMfx8fXKG6NcnvUw36CcZXNd9bnF1fz3CfCImABxlYc1i91Z7rvqzCxOa
38z0HLhn7JYAzqlolJUZKJnx5w5hzICiC4c2cpHJy8jxgFPF+9wU2DFmT47a6p4LIubZc7TwrZZb
ofa+Gkv8BX7WfAbPY0w9gvQlYSp6fLMl6s5uHO0JmmfvKX1aEBmuLObU8Bx5KQ9Q6pLUsWjQwurK
8nXB+GsjoBAJwaO2NXNTLAi6yzj8gOfauJkhtahoxTXC4FIh/2sE7VAbOeBjJKx8Vi6z7JcECu2g
dwHSjxKZw8Z/UqkHqsz8/VxzbKs83maOgK08Jtna+G4pvkYhBkz5keBTEfvX2/rTlbH1kztGpMRd
hMJQc399F47dXGUpYeF08PSKdu4zJA5fHEVqRMdJFahaBDnXQX+570Ba791WijU9mUDy8rYsNONO
c6KZnytnKuJWQkVzo30RL/EENmT/9BYd7e3bJjI8/ZGkX7ZC0l37HQL+Z5lhOBM1C6fL/wEkX6bv
wpFEzp13kwJrXbKkIoMnhHjjt8JcLqqxVYila6yNrdfK9FHDdH1/JynbZzi3QkLHQugYsRF5/BA7
kuZ8TT9LWKb9qge+c8IRq5cuTml+6AoZKftmKzPtPMVI3DlaysRBYAeIHGblUgi1OH68yydRrQ/s
71TbRz4xmK5QFgd2PI/Vv9IzPzZXhgcqGMxd/1qORfr07mg/31MUJe2Q0GOrMkiLTgQbeSg1PCFQ
VKY7j6X45bs/fWTyu1wDRA97ymxYj2KVA6PoKXpTJRN5e15ZFG+tlWaCyzMcGZEIwivSII81WQwX
Ts42iYD8NlcJw3pNClZ5lNGS8GksL3SG265V/+Mw9btq5HjoCT4CBm2SRkNGQpoiRc9pMCFt9NH+
QcrTjY6FOZQCccHnsVyr1c6uFLwRETjLCiLOH/TpnnS08cwghG2FkHPVBMMLrPUlR2MgOsWMbznA
BTCVgH1vNRGs6bh6ZcZg9XNT9crvTA0G9QHMtNrY06syZADjEcQOql4fYLj+pd+62Y04qhT0mJSM
i3pSRa/r06sK66Els8+AUN+nJcG9lXcLMxR87qEM4Cse6fYGLPhOk3iVjJCXwM34tI3y08jvCJVH
92UkjDgzmQUrmFhApkZ23vWyCMF9M4a6j0iQS/uOyRbc7Zrqj0pbtb0ISD3HtAbVtNM7ri72P5QW
xafBWnWHybOnD37S4Y5ZLBC/KRQlJp7yrP6ckPM/6XP2pD8dYQ4Px/YFI12hUD4HJ/vUb5rp+qgC
XjvtVuaztIcjHXoiTkLGzmnPmyskJ9NcSC69WVraPuqQb8QrwykiSbhtF6Z9OfGb31bTJMD3Yj1U
I4dJ/vcqGPi8c5pl9PwngHnWjFpG43/Uce9DIpjqgQ4GpUZeYu0T6rUb4+dem/FH7jcTQZlmkvuh
dlBl21RcTgaqTgpRJflepUmFEmDvHBFoU+3WZxeknkMKIYIBmrqgAfrwsCyVuy/GlYrSyN5mlopa
QA3a1A443eYwxuEy6UL5PcA6ADJChy9EYeQ2XBwRGJpG8Qas8KQGYf/bKf6qSDsH/lDvSPIwTmQ6
T6KvLcibyfBLsmR1MJdIOY5GQONwhtoh6nYW2CWNhX27ZL0sGuMN8ecaE9+8JYP6ffsJksOhD01z
SeZbf+kEqZaGVCXInct1FpbQyFwpjg5f602NHH6ecPliG8VT8XGFGa9Yu0lEFmww8wkiJy132KZz
PP6Br03SCHOdc1uLeHUW8QfoFKFayBK2b6IffBS2YScHYWCA34G0wXBiIo71lxluZo/yHCK5iPkL
OAAEXnMZn3OYVvdVllbAO7FFkYEKDLAQyqmtsG0fj/qknfehmXfSMmqoU1oBsfGUowpwdJ+gAHWi
tUolIdZB3iNOnSBgmhD9f87ugUZzm+QvYLPU9hR4Sqh1qEqMWaIwjy/7Z1V+1GxGEUit3n89JleR
wwxTODp7GFox4DF6gOs2RWQow/Tl0zosH+jKj436e45209Ng60Tn50Af1fx5vb6UcZ6HoPfzhd1c
aIr5TGYDCFFpf7DquB1eVGORn/gYss/TwexFBOW69W/Rj55mjSN0plZ+UZXUBxt/YmSVGQvJyM68
2yN+pkGZQTmOFgeVwbOXsV0UShuRKaRJa9E3c1sjKJKR7PeE85BUt6WW9Nq8rDLJgXaznvOB0uUH
esSnFAWsf430c3KR9V0d5GHztj4VjhpR0yQPgio4b3FiHV3H3eCvzxzuZaZAdJsmkX6UvwleKwn4
MXbjLYET7XdyrZcXOKzraENKrO4uLWxsHPm+pJne1tUT2Q7FJ5xSmvE3Xc0wWKF8I0gX2YV+Tkrd
mOqIr1SR3JlBN3aMZ+5AIEvzVj0FXWgls70SHpS1GrBhPWf3hy+zAeyqOBTyhL4puAOewFdWNU7f
6RspaGoNnLk+70E9yByrHuao00DFle/+9g6YQGs8WsoLxZn93C6EUOmMa1f6fTjVUvqvWZ/KA6PH
In8+XeYdjBmDbuYgGcXjslcpxyeZa/F8Jl43uQKSNOmTGQhodtiQ4L/st2ELDx+BKz7OIhy3HTEN
MOZslw8RnxiAbrPb+TB6kzcoGboXw3GLXgM0bGbOUyqexabe7jTyBD6VMUHrPoOG5kz+cSPhggwd
ZMUSuN32pRgAz+tyOLUQeVLRbLVkdz2yJ21gmnkcAbS0VTYc6idv8mmi+8+NK/NIB5kzjcltuys0
okLUHguDfWdGImB6e/pqvVBdaNYpxmi7Sr1J08kFh852cbaD/tfOHIRad2nWmIYAJqtz5W0CTztx
sXyiChgb09c92XrdiaDvKs6XrsRKSJ+y3lpsr/mNdZe2j/Dq9q3FczhQvil/Wj2lZVDNnGpPuiTb
pEjTykpJEhZ7cJv2Dl1obvi+kwGqimcgWoFi1HL95JhwNKRQAiEiY0m6RwimCFm77jK6qE2Grp9B
pAN2fOGGmJInikXSIdHdwqq1KHaQJEHObs2YkQ+xRXAxye86nyDPc4YKkTmkSZokdm6LIqFs3uFn
R3s2TJuKIugceQY12kHlA2s6sGbPSVDdL/rZuTxGODIhShc6LFrN1yvLpMqCgiU/hR/fYAInAOcg
q6vvJuaBs0DDs0TVev6cYWnkbJnMUxZQFDteU57LNOU9oQMLIF9OjHjdooGMo5TpmiA6m4ucO4Gg
tr4GFIDK4QaxHYkJeEUqRtmZsbJFAB96S2aVKeA38u/4BWSTjkHMW6mOWpZUf7O2F94R+nONB3uJ
Hp5E/U+t451s2udDyjScvWxE93lPth0B+r/jigFjedYfOH/ca7JpJwhiw5B/5QnDLK9v2wWH613/
r/txdAWKHkU7u1wNrHhyg0A1kVWLcaEmmJJEBh1dzs76Qm6ysBgWiccdEK9lHneOUT+FrCC9McZk
Fp2fZRi32vSYIutcVA0/oWvK/LW5PU2mrtYMIYeSNxQFMufNjvTY4OyDR/fzZP6Ep68WBXE4P+WN
PuaPCoQVmVPGbfs9wDLejTBM0gAsK7z2VoUaGKB6Ok78B+rNQX6lsZgpRDcwxczBRoyFtiGOe7jb
xvDm5CRlEtvbG70aC+KO3FVu9w6hO/1dIPj9HOn3jSa0uP7nED++gisCqdIrMyPgE+lZbqN8B9hT
QjQaxiGoj18IpuNO+4HAp+/Uiu4Po4bt3kjZiN8xMeNMCVsN8t4wLl0QRoSfx6c2+HIAxDX1XeD0
hSeQd7VqDVNJdKkV82kaU0XpXzB+TyTLIkg/XP8U/K7cDIT4eCaMnyDE5f7lySkx0igNMi9VDG1u
BSlAvvKu3uFp5J1WRlBbZRcHmMJGBuL9hJhXFG7FZWvo5MLnVGTof8k9vAxbZS3Ij2TCBmx4kRfh
SXdURc5tsUJnQtspIktgGEE6xAh3pXEdUEfNtRnS62AEXgLxWi+paOrKrAKnxhf1MiVD1b3wegQQ
OSbdDEcVglZ0u0DSeARLJJ7mCm2ULWnSewpcImyqk6TIkb/ns67e/kzxlLMZWQXaeFgo3C87FHCf
qCHPrSCguh0U8BVKo/AoP07Nf8dmJmZb4Yo4CjqZ9/xIlXbL0DLU3HbdmhwZ9vxwk6dJdm7kkNcu
T6uueRQPQTHUFjzux2cG9fclgb2MVabIWHZNCbUXh19oV6gfdj2msB06GsiegBRbl67S1Q6T2gAH
kOEJadcMIgN3LM+SUGPCsPs1ZVEnqjfYR1pizUxCpqvpbLa01toUZ8ebHEVeIfp1HXBlmPZF0hp3
8lQ/ENimP8vC4+drD6fEl0+YpHYx7WwuBu3DrIsYiZyQlQd/Qtnd7GLvNkxwx/rhOC5hSqcmE6dp
CVP0tH8IXx/9CADen3tVjL7XucwNebaTOKAwUWABDZ+VwKISD4krl4MH/nfUlw/cEXMt7mcfxzNk
7o4wuPGnRkpoxNU03ruLEgsNDHbf/odrZKoAqIFgxFOPG3Z0dRA4jGWvsSSu7l8goFQSKE870Krn
2CuIrJ08MBbfD/8WBHuAQ/dhe7crXq4OlYRMBCMT0Zvd4NUSg06rbhVMh6ODh/BxRMPRiaLKt/8B
H0yjfT/VTzdtxvZGhZBmSdr4XBExxGoz3Sy3noOkT4uEdBe/P9Q3Y/5+Sgr8yKIyY7b8LQOPFWcw
Ne44K16NYwQdEaJoanK4Zuos5TpRH2P22+L1TegsMwg9g8bn0OMSB31e0NKmihmeCzZegbcT4zYm
edgmv2zWoj/0MTAlvgfRIYY/qN4UbMX4sQi/wcSrhboRDkGNFEu/R+4jOLS5xMuVsxhatfW3kmAb
e8Xmw0+hkdMkEWgewaeFl4GvNhbOusxyQzypxiKfagioOEZFTWOzjs9cYMszAmB/fMkIJY1pMTLL
yJpDYDOmH7+VCmu9XgXdmlv/XHptvDaEk+QTzEtAne60IDGONS1h/U1OP9XeMTdF9ztsWEberi6H
cdwlKlpHhA/mTrJyxJIdNBE0LuhSDUuFhUV6aJRjOa44+5hSWI6mq36K8VSc3ke7feox+H+YiCls
7J+vtkM/S1bOC4gINMvto5wr9U8LYW2/WrK1Kq9qO7WGYnulNUEg3sqois/oFDzFxJPohl9V2vgO
g1yVo+JNIqGNV2BY271tezKz5ujJyGByVUplouL+Cf2kC6eC6U2V+Rt5I5jI/WM9K4xKMg6JRc4G
GAsLKADN72a4a3WE7Sqdwk1loaAS9bU2A+K+rT83RlYdKJFhTz9omn9kyVb5GPUevVqY2jcg+vo6
IdpZYYdkq7uvboHFfbZHHYI/CsLZ8614naW3FtHimEBzxNUSI8kdiTwIm/m3R1buDCEXTJaDuYMC
VRrsHrtjiLmSAi4TGM/TULYrIMl/RFeMvjQPkXT8543gBVejP3WCYUZbjfnJH9RdEtFN3rRAkaZ0
oC8jLg1MPhWDdbRRd5vCxgFELUQafm9yWaP3YBovdEm1/y85j14A1inRQjmHH3EmYfG3YHN39JO5
swcKsnfJFVlSWXOyjgNthI1DDcgXnkL7Mgk7GTq+8zo5G8GB9aaVyqP912cdOqXCUMbmjeK28l6L
Necw7Zjb1D4XtM023XEHgYcd4Pwa+P+jVW0MFYuqdPmeyX6l7/cvYASR9GvyinJrGU4q3ksCwONu
5fH11BwVIcwl63cQuDEd/2gQPC3CW+UunVzNcvZ6NZIjDE3WtisuucN5zXHR0Jp1LyfuWpGaF+G8
QMK8Fqpmz5XqYAVkNSnZqNoLANs5l38kXjCsBOh+uWXB7BLAZiBrHT0hsIHA+k7d//tY8AYU1ETp
u73iNMAPsEfGehOa2Z4NQ0nQj6c/JEc4YgobKrzHHRdmEDbxdMFTvDscxYl16hiaZlNxl2bbteIr
5hYR4qh+0e9zKON722Q57GMwq4vQolQXcEyQcNjaeaPz+6dJ5iL7IwzDaN3ef2JXH/20loFLQQ8q
US9E2vAfceE9M4UW/l3OBNEGu+Gv+cv6q//og1TzUMrkCuOJ/JUsCbMbD/feZBCL1Pgm/VhHM4CD
G9mTmMQ4FyL/1FjP4XlbkUc+HBAa4+09RdQw5beIkq+M01wwBcfn8uipza3CiOhWkrDTg9Kd9Jym
Ynzvh1/NMwkCONYQRyaeC0TUu0+4EraUtL2ft0tLRleI2B03BV2jwCDYptbXXaZkflGPkM1toSPS
k4I3+tOyaZBhaRNV+oNoVsKd270ppKgr+Aj3w5MSjAbt9vy5s2xA/4+1TOyD19vylZb9B+DCRb2c
Gpl8ZiYuvrfEiKBKOZM/xVwZQOGPK8n7j7QEv+v3Q/NzQsL2T9Wif+GwVrTF8Zd2R+mFsBYCpm1A
/UqdhkJ54ofKYmf6YG5gmZBr+1uQ7Aa+oqn/RdgIY/eUkagGUqDEvr3epEiYAuzobgkDJt0xm4LP
VgY4fo0F4VsRjlvHTGdTcHG4A2eRoYxUxkMMm6GJ4G5ipv5BwqQ8MYaCEIZ/glETaz7ou/T5vEQR
s54dNtlNmJpg/+f4xuu/QChHfcBH3QupMQMux46uzes4rdJpBF94aMoCsqUEIdjmKCKnwpE3Fa/7
X1OF++vmGvvFPrSRjYcO7+Uu6PEtApBf7yDhac/NHvvZaCOqjGYXNSGBhQI1yJTE288dLKDusul4
3Cbov6h1ILPjmsh+x0c13F4v6clV0bIS74mGjoaRXx+5wRd1VT+e4D+524NUg048PFGb14BiDQV3
2Nrf8vLrpXsC8iB5akTBGFzEchJ+5D6ODrBs3sK9kRQi9tpOfUtIoeqdFD5/GUcJxKoZUcTjtvQz
37KJ6UlypMFgVYGzAYBu4GoepiB0E2dw6hr67cIiz7WPtcGJ+8/qXAwqudEYSc+USOy9Nf9qa6a4
I2Tvm9n8X4+YhS0kWTsf5yzHlOr7iNbNQ5IC6ArajSfMjwpWhAjNvF0/qPx/DZbCeOR6FdtfXKx5
KUv8PW09eI7UfNF6Aw5MZ9pqU1UeC9zs/R2JhKrd6e2orW8KYWEUaz5T78KQJYfL4C7F5JnVYgAp
AEPZ6xv5LOATJd9FbuI0RWZCY3P1iaP/PiFYTL/Qfl08btx2STPeyDzvF8lBzbiF5hlFxK7PD4vR
Jl4gwiQ9slS1o3xcdMnya6RoPib1b7D2brj8ntPo1DRBsjioWUD9D8dR0pN5u99g0TziuC5CnvPp
nyE8MAGDasSFJyv/oZHZraBZ/Sj33SLa4y3kumTwMiINDQyoejG6C3gt8D4KyUnNd9ZHdgrpKni9
UlEO5AP5eW7rOIlYidQLfCbQOS3Zz99c6JnTCZyGKmJ+oiz6VJAURKU1zjBWQEcD0fVy233ydr1N
S3SQ1/AofvKKRWoNZxlBudTGpSRKP7c8Sjp+iu95vZGImlJjUDb7++llpG4LTmkeYXpQrAfmSE0n
WBZbR5AAozJu9/aIIuQg0hwcW6I//Ooqe1U37J/9DD2q46mCiBmeVynUZXsZ7fVCFYQyIMC7WnsT
AJVWi8GovFk1OImitg03xxC87Ggp6wj1G7s5L60xzCgYJaR7OkXhaHjctvk99tPyJEmng6thMhYh
Co+6v/KOb0b1tt8rEhZJmpskvSwVpr/RvPHnvRNGNSVuY/S/yIYGZy2Yki0x8FygMrvF+3V2DmQN
DQeTtxm6wQLi7CLMXU0Q+/R3Sv07R9rTq5dO6CQKqUuswltE6tBEWvNmRUhzjf5uhox1Ze1dCsfI
VIcHCgJ3Qy61uRyOTd2yb/70zdbzAZw+vBCrqz9+AXedV+tzROEYoCHSjwBBmQGUA0YmodPbirsA
JrBpDAX8nF61Enn9R9/pR1QeRw8cwtlkg88XF6e81wnLLeYk7UcGvgH0oL5sJUrc8205JFwiUbtL
lO9eZAmykbWLyeEeObXwEFOZcS0eCiSNo1xDl8No/HJAIouSrm4T5LK8B06yLmX3n7iQHScE0V29
/mCkKFUXZVAQhnVIk0MvMJbNAOP6WTD+NEQ11P6sS1OF3hXCeHvmIHI6YuvfxzINGtAZvHz77fyt
0OwbH1qd2EdCak7k7Ow5LfLBeBPM8vMLVKbTjs7DI5/byG0q7NUM9K7v3JhMHCsaCMsm98mabiHh
Orr+BvkgPICoJqJBeexZ3/IRrNRxE4JdAFjpIDaxqkkIh//HnCYkE2D14Y6u1/HVMoWjTa9ZEVVh
ZfB6tcWXbeGxqI0LvvOvY1GlgkP24GWBekyC71tBz0iIxd2920MZcN3OOqN5qtDdV2OXsx3n9kf3
J/IkWLmxnbVgOpv+9t5P+G8AfglWOCDWbQXNdYE1waP3q8992vCQi2AcVsdA7eMj4EH+ogLyf5oE
wpeNVpt2KVxIxcCXLL5k1q2zLUQ07j3hmn9NS2alsh1P3vKhfBQpoTTAPwrbKbmd1qHwtvW4VyJS
lsvKJfcBA8q6Ls3YyjPA0VKNTwqDorEPuxk6qdt6rDDxe7TFJMJWUf5SAog9ZVMnx/KOv7iv8OSI
5VD/uqXUxGlZ5WfjgW0UCiBS/v7CszXBhJKt6LR0bpkorm6QgZT740nbFZi3ic2yYcGzshpaaGzA
dgE6miWGfECLPYq78bOwuFOfSCZ9oTzva2DENCZlANttwOyzeTfzAS85CihUdyCHRS3PCD8Bh768
T4wvpvli+daq3dwAjY0jWFpIkPKPr5VplyKvXzEkOIAYQ8pGfFEjjb+migjdwu7qUUCWiyI5b/Nx
Z+rSVuZbaZHRFrD2m6gpoX+lnLKS4aj6N6sUzVWBgMQ5og3AVO7BwfgUjh7CfZ9QeJ9X2ATkPdJO
4QTeYXEHdb6pRQX5E/JJONnpwZCUXTboUIy1wUcaUmusiKjL3JfU1tipINfMTVOzVz8i2maOJYcw
3HueOvTAYY8TiHPVue62qUbF/3zwRUmdDmRAxTullT1FaoXtTlYEXhQuu6Iw1qGL7vMgophTyy2X
F2PU78xc4vO3EAhsmLwNxOjZrwQwzktrl86E1dQhLpEQrlO2W2H1WWES9oJc8F47feby7LK2DhqU
c6wVskMPigeDkT1Mqhw187K9eK1XM3phMHnPV9FFMYW99zHyLdVpR6ZId9cZu8aC5sT3odrnEebG
9/+ZUu+IElmZU+qXBzIZUC0ohhTUk1+zsre8KFtC3iNPLXFjKo3QB33OxwIIKAl5gimz/rQeq00o
v8tDQ7JMUeGTRHBxuFX5qf4XAtFjcZD9r++rvXRX4twccE9pbe4G1fPefw93SL9S2HoSaY0bySsj
icWCrn1+cmnHHU6/srJEXcEylc8wSoDswdv5ur+/0UqjHt28RdUv7faS4RR6nKpQY/9vx+cv7dOb
Fa7PDfNTsBuAsV7E5IsfI9H2KD/tu868KKeaoc0ZaAwEtM4pNGMlsH6pjZnfYYumceCRXmqH20rl
c/Q1iM/IvXrXvGY6ACt3XpEnMFXuodleRvLB22s0jYdup6Dw3/Ry67Inj1UvEuBQyC5sT/eX8fgp
L3XBfpDaLDz4gDPpeHwcWYNFW/LeKd7ZTamKew8PCiHPyJU2LTpqIyvV9p7ldpsYLBUwWLjOMR1j
P/JHpdzAFYnx4vPs7kZdPkl+X5GN7brVAVi93BvXaHS7wfSfpX5N8GTb4/XIo3CMHbs1aaTkiMlO
AuYcw5I27YqZOoeaeFfp5if+j2Mxq3ur7s12ww6Djby+MlEQ7xkCrn8yxMaFPv2Yv2gpxNRow6TY
CaZt+U6VVSt6j7+7AIPezFTugoUkD/Lb2uFioNxKTinUP1vUPPGfyXjx/5zdk0UhgMTdXVAwCpjX
Bf3US6Eg0ROYbYPjk3IKnwFGRw7mji8Ez64NTiLwqV7+5hwz3ne83UDZXJfbd/UBOrkNBYO95Tc3
k+bO87j8jj+2BzrMRqjAxezt18yM9VfoYCcZnSNHbHGa/itpHLHO5REgNtrYqQSyZP95wQMZEIeN
aRbiJtb9VRgmzcl2ziwo93afIGNG+y+F4cky5d93785BfU1TAq9EGcEbPylspO+P+aTpOazzZqRo
eSEsRdYGzEvovzr3bD8hjjGg5O5vUVczo3xWLgiv5GcVSVS3etoJEnMDJdlx2tx+1qUI9RpWVQHp
W7rtwQ6WHqZbqyAn5YOKMylr5JYfdFg6EiK7ZZqnhOauR65soG1tW0CYuID60Y3NJCFxeEyVWvx0
oe7kYt5HUxlsMl3GY3lcjBv3XxL5HQK2RwVeGzGvJLfHaRqSnV6HbVyL7h/Njo+nCdd7GHH3Fdc3
+ovfu17lI5kV4qEVDL8NFFyFrj8Km5n0mPbzILqsdacDNhmP8QB/LeGR1Mj3nrBeqXMfeF+MuLLi
9F1oPl0HpgeEeURKDgVAf9Yp4+63JyHcj4nNs0cKVWjv9DsERrOQO+biEUaeJ3s5b9+JyGRet5N3
lNLv29c+UPpv3bQ+mQfTsjI9Y+/Rt8txVq3LyLg/I0zOCQ3Iek9Bg8QD0fvCd9d1qLa+jwRD6h1W
uCHjj/+9fmYGLL+xz0ng2iIFm3R2XAzURCB+IDwer8ohAgyyUIHJNwWvGq0j8nDYMi6YrugjFqwI
HMMCuY9VG1opVkAHmoL3eC5KroFE2xKJs0X/4ncw3km3eE/Riag81r1i90YGZGn3qhCneYGiV0pU
2/gH3lC7E3xOUugDe2U5x9Wclh9mB0aZuPlZcu5h5t/xkCE6pIdcbT87TjEublhyIWd+p8Umo1Q5
8sRhpoYsQB2qv/ZIdlQvf/yhP8r8LgdcW4UZVu3ajx0epoNxtvegg2sz+sqDXRJIob3jYELW1Pmi
+aID7A6LAPX1GxTBeVTFcOSUM1fhWMjTPxr8Jb3uamQg+2ttAB1SwY84COXP8YtbCwTlAeOmCvF4
YBrEi6oXBFoGxTnt40Noy6SNZ3BvFLgqmwtbHFdGugX48xlEYWIlmERlawONbfonbsJNzGy5Z9VG
fFe1e4cNKigd0EYnCK1XsLPRwVrH10OYdIqzd0qKREK9PqsJlaF8NgV/a4Ak2fyhFawkn9jth/fa
rLqHn2N5ncE4mKoXZ/fsuDzYNEztlIOemyfuvh2KKaoSbUEg7xD8FcofSv/5Y/3ygi4zvhU2uPFD
JL/8zlcK8QWTJib+mByRDldULkk8AKc81Q5xZ5pM/Z71DlUC90O+m3w5fgXAQUd9mKavmnxEcOqW
dsvDjyPb396aSWTk9zYVyJaNvoKYsJSk1dwN3AaTrSya6nSo6NqLYNkBmHVM3yEX0oH4ncmsnspQ
jacz39CwxQq/YopG5SiHjKbkb5UiT89xTpJ1lj9I0J6hVCkaH3fC54isljJalaDegHIcImdOmIFt
5aWLrcthQYGvYEpd6qk1cxY2NUBgssvA/PR8+d5SOrSRafsRvOl/vIfrhjHxvXK0tO3jnMeULfXg
HSvRXszKKn0qoKkxqwUua8vO9c03ckK3U1AzprjxARC8qF+SYasKxPc4mUYb0cB+5j9nVDAx51wm
Nw3V5BtCgVYBzPwZVcMsAGbMSid0XtTwjwWZtNl+GQPXUNkkMjYYah+1RgRalinPH8pELB6nLMd3
MdlMbtsp5XLI2KZABE0he81mfTv/ksuYbpUhvjXUcLtAB2E9GluM8izmdDNZBbECP/rAwtJIjfOw
NP6SVyD1cMVjUdktZshKH9L+zHJAxnQh9veGfl/y8N/+3XtrSDbALAYHt6N4n88Eb6vQnmSTz3ft
q5pYqyaVKFk88gmCM7rzMydjNmz8cNxh6O5MOcU2nBNCLa6IERw3BF4Clgxy1NVhH56P/TOfGVmw
kj7tnCLLirx5/yO1Y33z2n9EBEvldtJs1Y9rPmil943WPRouQ36wUIkHkSk77tg2Ipy2FTcpCHn2
jGXVOPgolaLiUzXeG7KFUXV/rYTtr38hYewVcXQSTfBzGn5HwxWQSMQ1F6ldABmq97C8rJJNGMRu
p2oFW9NmMTuLDftCajUSGOmNVdhe5lmZsnao99qCDQBC3Foz9mwFDmpYTokTZNnzT4X0zt7P8YhJ
RdNgSeqPEoh7S11/TTSgA/LBNFilSs4irrRcV4KY7ojAjw9M5RhyE77tA7P4IBug7AqKSxNSJRJ6
yD1TRpZZoBW9VN5XR1SuDax4r61mFln9TrL3HkHiGY4OcyRD5BEEd1DzuuoVQhlX8pp/d8GuXroe
WkWL2+5nYctvlQXBXicHD3uMMZH6XrV+8LoYLoDGuOrV39VXiCM2dJSZJxd5GnXoAPP+1yje6huj
AuToUcCpZwpJksQd1ojFmgwysuRU/VU+eIzkXQ2Dhh50YwK2q+Wk1t382kPP0U7qEJB4YpuJtIEa
QJsLiZQGqYmtnSNSPI7z+u7UGXytkqi+YXyyna3bC7s1hn5e5aHEw2m2fMVWDkodPchjSqN0tfVD
EiKrhEGDJELx+P9J4dSq1TTYIOMHXqP1jv4lgPCJs2LnMMkDYYVa0vevZQBiadRtVX3ZOZNDCBvF
BqDdQ+BgvoMs5/jnOcCc3ydVN8RpcV6LGC2TujB6AosbIJdGs8+lMX2Ll74txmP/t0B5yUu0GPQq
2hvn+OcgAvs0wYHJk4cd/YsWws8/tgaTTNIHjVGermuvf1XAKFAE2z/QwIONmEY8O5qNEvO9icYU
xtrO0UGEvuURkWAYITTCT4MsBvs0FhLzOVM/0GZyKsgUOROvwqmcQoDj3BrB+OPhpHhB4cKysHNe
5VsVzRCT2gNFyNI2HokA+pFsy4OpGFmdI8CafV/Bk4tdKMitFfvczNTID3zvDAGWokpeDPwUi/5u
mZ1pNpcqU3Kfk6wTd6QoYLwTgFXuC67+cL6x7Cw9n6hQwLkr0yeFF77+8M7duLxl+cXaqCfRsUn3
VmbGa1v/flF6Wy3YVrfxKk6f4JujCVSE9j5laAoQrytkjKY2PJjKTDJyFi/B96pyl6Goddshz2ZR
H6hcSbyicSTIEJ5HmD3Oiv0zZCnTuV4+hYiYhkOpo3ac0D/pPROKqhEjMQohGQ9s80kqlby2VfBn
XE7pxt5VZuMfzcXYgBnrjbrYceQXmRVzGQozSbNlhqPN5KLoK6tcKnDvkDIqgDMM4JNORSUI63vt
INE4x3gNaeTiTiYgQokYa8YvWWoiaWH92Sw2FIQmrO+mCLHTtftTmv8j0CMzwryJYg/G4HlHTx32
+yHnc40e5rLE8+ibQxRUFP5XFgQC5PD6FJ5cmKu1u7rAB1yFfvYHwSxqr0q9WIR250rn2/SCWpuK
KzNlts01bKWQ8g/c8IrOxoJMkiIQ78Zavg0RaYXwdMbwxr+wld7nGTBb0jc5ScX8D4UgHEV8MGMl
ju/Bh7H+bgBTmsnc6sgH3EM66boCr9SP9OFhwQ8MbYqOlqaMVlOGISlQd9UZzygnQNEB+5KGgeI9
Zv0SrsSwuaTfcY3ikdIQoXYm9rDFQ/AsPxMT0G/qaAWPXwtDK7XrJ15EzhKyKIeVPAs82qU/JlTd
o4zs1NISHdcSWuVrUSnxl+clrWkhv0edJOI/fi3EgTdUODU6YMJwRKWyOVRmgEPIzuSQEyMjzqvT
oB+PNTRZSuRDccKHA20gUsEPTxiOItQqAFanm5BbOAlt5aIkBRTaWODRt8VyNBH53aZZCPdZfRij
NMG1TOqKY5ne07LV6ARPGFft7cx63TAqtAEw/pSvDcZMlAik/Yyhq6PPeGFD7T4ReMBQlCVdlIzO
1sUcCZxts4CIecSCmWdbnKD98PKgV5W6HKrqQRHi3eLoHsNPWFUalMcVz4E8MoAQeFfPmOD50qGk
5RYKYCw+qQI3bQEcUSk6JMjm4HM9nPd5YhK137LasUS2nLGI6EczxHisf2TqTObJp/2mbZub2diL
O0GSQm6ymi4bH30dzKwFsYY4mpNF6tsme8B6M8BPl6Qt+h8GYJrhiLB3Fw0G8OXlsVrUVCyElsk4
lVlsmqG82T5lZfc9A5lQKzWDTKWIA4fB472bThHxhjbkg7sHLrxCKNoPz443or8divtT9AZ50Nge
391f3iCA8hk6FmPegAmENwgFz6SufzObjBrGqAeAQ/sfSuusO4kOOx2/TVb2bfZzfDDHhUd7tLEc
8FpBZBLXhLwgQPw2FodwrQvM/PLQ2BAKhCWrQhqTH3myMAYjXdNyefHwdbfLPr0CV7dE0jz8KbG9
2Ipj/dZezdQjphy77hMV5Y0/5keMBaGYHSfhiAK9yr61MMuCgaCClU50zKXH+b27d7fhAPEMMCic
01jdXB+r+x8QSnokTb4qHmY58wnhESajI1N3main7q/IWOLMFF4R626FqInA8tCtZiIeBVXQRk67
rIZMzjlgOTT9/Q3KM67PW/URn9GR0G7UIuQfCgayZqOpJ1PttMBTuWXI6JpSo+txqrK1nvkOqz/2
xczuc1xrOkCZLI5cq5bpTrMXnsFT5RI62fY9l5C/fS5Oc/K2VMBXl8iCmyHRsiTTUNtsD8GdISes
lGS9PbRUT+C7ekAGzbVA5DOF2Uw0+fWY47hchA80bLYFGDFz/SbnEntjU1YaQKeOuyD0hVgJ0GP8
Jrbo5mEeTvI5PMwOwMwY+z2MdlLU3p3hk4pwI9RUVAiYhqKugLyne9zCeEciO94B9/xCaXrPAWZ5
FuTbqPsmCmr9MDb8JEpfq0K1eu53ZK68AQdibRv36ininK5Eg7NUgBrPTh74e3/wlAHpcjEITMxx
p4+i/hT8KJ/sSZvdgMH3JA0FahokNh70ala2/eDtLBUK++zwbq/TW303FgQFYWQbuYkZyi1V+74Y
uKdj14FQX+1MdX/Q28KoEBWtwNrvJFvLzA1ef9spdXcQpHevje+FOBw+fbzDA/puu3ev1xmUStES
YDNcOEFNMbS0Z4xCZ6nUvcgCu+6SYaIGtHLDYcZaFnzLCP1T0fMIUWkGf4G/eo/dxXb+lb2lXwFg
9LGChfBrdWf61oWLMo1SzIIs7rMLr7GaxrYKHz5Gk8pfO+Bk/Jw4kxCJR5PWJj0rGizSYR1BNQWf
xUpdCX6OLx5iwF58XHpK9CPReqXlVOl5y/4qQYMpBc6ImLij3Micw7jnYJxKcf/L8mmfODteP4QP
u3wnxCiDbRsPKhRKXLEKPDP8NCIu6qIAYXncFzaUF4M3zX0Cmy0C8px+RloXlUvs/eZgeByvta6L
2Lfjcfu3h13132yhCbAiap9vBJlwrpadqX6G48Aho6kxwMRzhBubZWq6QDhMzRM01X7CY1ichfXK
jB+swzqIYQKUMbfqWEYtNFrWKXxsoqGeptwKq2IWfh2Oc/iycaz0TodQcaZieycH5kEwpZ4lxQ4k
FhhKTLVvUvE/b0ITAchCG2xYQkBj9pr6fgBiedYjqHDXHZ1J3SOJgL+cVp1jRTPD4Gz1LdH8rhCw
dRFxJjEbo3VPx2MVyv9cpyCP56a+mCVMt/Lf6+j5f4ePKQK29hEdh8Bdi2ckd7HsyZnsV43NpZ4a
fMP1dNQZ943NtZPL9wiWskHuXbI+WDUVrdy2x3xZ5jbeqr/fktQDpBSP9EGY/Hj4kc2SK+jmJ8kX
g/wU6aakCJk2/YYUKrI6NmSt7aAxWx5eP8Q53XCzFk1z46R7qPxBOxoQOvvY0NbrBdtnkCEnCqP9
nt+DepTDhA34EpPbPb1Ci1xH/ChGYcPZSY8iy28UoyoXTJLGLZD4JtVEPw2MGX3+fmW6AbcVHn3e
CfJUZye39oerLa1mf+NPYBZCclcOi9d8r7p/36jye2VEsTschxE8f+hm6dnAEMKnjYMYBrbRm95C
rJFOMXISmuoDLUbeIliKv1LeY+RB/I5MRZQdmBz7cr+6S7h+redy1ZakdBj2lSJK58Wsvhdv5jCQ
gDlC5VQtU7rfaD4rLa1rpTHFLrLbKLbLpA9iONvLGFGfN9zhY9Lgm9qE5ROgZiFYjdISJPWHyCRb
mjHQabuTXvm5/P5XIQEqE/ifxLhLe3RukBxAw/ZPAFbvgryxbOoz39kWiTvFwGugEG1y3nSt+C/c
m1KI124FkuMiKnORh+NwHa6cAwEydK10jLkTYiDEEo6wZ0PbsWB9tO7oRfLp3VTUNsTUjvx5Jzc3
bm1Uf7Io0IhdxgbN8C/0/RC01kXtYA/EDkK5x+vYWv3jP5Gr66et6bHcxcSdNSLqXGlMF4QgfT1H
LRsesOh5lggeocCsC54d9+7ee+lii3PZZQLvHrCCE055XxO/RY/N9FrWx/QldfZu9ncn53+uA2d8
8NmREnMijJJtrVc4Dh5ZFE+x5dxTnF0VWCkx1bOVY36Fa1OQtsr0rvoTqUxPHzll3vU8iGGjSuS/
hO4HEczkhE5LnN+2MZPEyzwKCjMqGk/ao0koGvF5j3gT+alLFminFuXVmiRwsT3q0HlQQUkAuRDm
iyGjUkB7RBpu5yFmOQJnh8DEcvdZTb7IZEIoTC+mpMBx0JDor6XE4XKAYNx+z9oi/AitW3L2+5TN
1DaEUUdDQc5w/QJ3Ajm8dIhhv553nK4nmK0IqojtikH1mUiOxafFDH/T3O2iO8vxWMcDPn9LV/bx
ICnZyw2cokL0uVio0vXc1A7jEEssn++mrL1Y4ltZgmwG0M582/zZcVvoXNroBSUrqyhwZJiix/IC
wtoiUEJAMztgGz3tT6YRbKWXqXZHqi5/1DF6FqWYdh/4udS49hgWy3kf82ktgCKTykYbxwkmD8hB
9Cc5Z8uiIz3PecZvPV4mYarzNgWoWJQHPzAhVwHGuLsfhfKppcCVC7nhute+LNMDDCs3MPBJhTX+
CIiuwqzSRZhTNZ+KeHDBcqFgvwN9IjWoQW3lh3umLALtE0Qhms6txDYyKvNQVYrRMHyDK4IVeyDv
j5icc+OwV+7t7myYfiOYvdmsXjtJTh9BpUBmOw5W8rPsOaO9dYd25xkjWWdcX+k0RkD0LAGTsORx
J3oOauVrjVjZ+yEVNRdlUtxqb2tO2UONqudfW+p1rFbZ57EOWZgpOXEdgisJAOANV7xHFzXWpUOU
Arg4VOLKYeszmBUqZ5eSURo8n01qwO2uFfu4YjidHNWjUPcCEDCBsDmThzmol3G3i06sV9FHddUV
lJDxfchf6MGe+T+cxuAVlh90bcsL2dof/22l1HV6TRKaT5mDr9a90+ak1AcaRk7f+irTSsVD9ETZ
IyWBbF/dB9xVKTCZRhXx1VCB723m5hExzuaWknU+0n1d2EipAKR+48ytTHTrrASe8t21sMtF79gu
abN/HpYbIAIcPvQqZqfFgY2YnlAofxcBVvt3gEqiAJmsQ7EXB0QIkJHccriVcYsBly8U7lLj4/zD
Ima+ZgWt+hs9J83nLYaosT3VpFbEm0x+pbfg55kfusTMBxaL96Dz/Pr5N1ou0yj6My1SUFuCdISD
tFZC+jfdGcUA0e6g6MBVCI42wGX3C1R7Zd6amyNsRUTQrg6ZZiAWv8944z5e7ifO3ANIFzoNAp8L
WCTxtjau7ilzhMwbwFozxLbJbKfNdneR048W9HK0JsTIf7SmPd63NxXYsd8coP3hHJmCAZhKnlvA
rvJ72cfAv7XOL8XjxZaCNe61ltF5yMLx51FsUXzBfywnAkoYf49LhqvkocOz7F6R5b/tFsifTh2y
OaLvbnKTURDHLP6KCtPiA9rWnJzrE2H0pd/WPBOkbgnbUXUixS79HVsocEWQh/I3woxR+c4P3Sw/
fzkGmn+1VuFNvcUWGOxc+wJMvdkOmqZzNR6Sw7AiT/THfQf+g+J9R1MKL87dtpdbQcoIuRkcu6dV
wszt+8qZOJTQ/wf1INvP5smZe80yInlLTGXNQTzzVUXEGu83rL9Oz6N9fYBguVREIcwIPBi6rQd8
AxUfaGcUKA3CH6hfX7lDslTcd/IOvEn6X0uqbITeqhrQjWkOA1FzGhfB+X5qRmCowCnS3DXiWmsZ
7jHpTjVV/C5XiOE0o95lwS8a1G8QZ23pQKFQ0G08LQQ7CPxF0cnXZxnRnSVKVlnvH1LeH/5Xesik
hA8MCjSecQvlzT7ZZdxK8cz1TF1Qjduz9vfzZKv5ucE4FYeLGSiBCPRUWlV4O4epe9AdPF8SR3fA
Ju3weN61fYdZUbpIzZQLFs0fVS7DuT9Jv9c33TazPvi79FQinC6KGBqLZEVFCzRwwQTHJ6zhelZ6
lOxwSOvK/NitoUcLSC9HhGGnSDYYzHmJQIuBhDFQjMQ4zvaDEVkHcImAM/VYRFtPHYQmpdpNpuw3
UKfljO5+oMwpzJCrPcK7+iXtVUIamYifV6ozXaA4p59JnauQCqsruov6PVLT2zjGVWESedR3gy2v
pVdQBU9LtnK/zpbSsmK4PX7xznUM7OFJ5FFKYO7Fi5VgR9MXleHw7BAYGAEKMjzsm1Z7kS4vMB4Y
zWXdkDvOzWz5nhhcX6zC2ZOojq76J503o/NXjTROuBBNDD0HUjUnmdlUeuehFEbaWWf0tQEfGFks
Vs8LYFBslnXwjPZS8aqevqFsg0EexYRYbEaHpCuWcPIwCTEyrwT+6WBpY7/IeUnqpuEUxp2TSvBY
Uorh70IYSJL4nNLL/Rjg7Cjg8hHwoiqPWiJsj899uXH26JIqYgZJOhJsQAqSCg09i1P03IFg9SWW
fz5/yvXnSBXYWJizuYZ+pGXfQyyOGS+g7VJsSCrvzhgvuwMFirugJIecEg8o4FbmyAE4/XH19Kpw
1NOkN2K1wb2coOYUo7/UwYtFNATOL+57jur4lphxkj3elCihbjF502lqD045nTfwWfargprA6V+s
T43VVDD83HjbyJKt1jSyEx59FtVD5FxBz86VHVM33Fzm9soiiiY2Y2EhUXU19uRcU+NmYBozkvOj
VbF76ahY5878dub1mDPZpI96sDkCyxqN7dIRJdXDgqA3SFy8ftTIG4N3Jt8uoNdLyBKRp2Uzn/St
4vpcLM9gVQk5/xadT1IMdhHT3T/BF1GOsWn+7fsX32U4txUKEG2ueiAQM+/MWsqgFJcEo4uPD2hA
fJky1HL3z5IemL42VqTwFFCoD7zIEkzkxiow/Ts3hHSQoJGq9fKS5eF1puziH3OoQ+RkqCwNBqZe
BjK+t/4E5Yhy4y6NgkgezI0ucs2n8aur/L2F4Yhscql44NgqDMGezfnYRWTjrYnAcCHH19DROWz6
l3/IAZ7TkVrlRkbv7nJg8ienjcHw9jJ+k0X6UAuocIYZNy2lAxR+y4Zj25Tc85a6DzkC+u8fIQn0
GsAq2ryl30RsBsE3r5cdYh2qWXZ/A4RDoSUSipNor2uBti0G2fncs9aHRuYSjci+rFRjgk2VtgMt
NZsak1YTx+zXcvlprI6SHwLUH4g0cbgP+x1ppM+Gl+4U/flyTcvsw3Q9nn7Ud85AoAuW2kMNoEud
ZopAPoMIKZxn8aKpbAeE9ZQyTgtZqCmgUwgURPLF85GbPVyDUFMaYA5yxqzlGgU5Mhcl8vzpDUu/
DTOFL84ZaMk9aGXZelQQx0KT6pAvAJIHFuMaStPqR2x/rXdtedWyDuKe/yniR5ROZ4PLwdSCUM8v
jY37a+poiY6KdGJLKW8hmOSpK1FCiwfT+bEhkLs9EmiPHHVy4sCj3lmXzdJa0SH79eRP+RI9PuZX
O5VCqXhnzoLwWhtWD9N2GH6AP+rpnoYLdeea563K1N1ms0ZYFn4NAbvbcHkqFUh2c2+SfksqPmEz
rWRYGm1mxuHCMHPlD6KWzovejnLkMHGlIUS38GhMqMyRPyDHLQOwH+6b64rBRJmnBajqliO+Zdzs
iceboOIJriGxj0FzG6JsjeaWB3HZ9mmCjgffkjEjxCR4zycfFlBN4tga52kjlFRWAKIfJ4xN813R
5BCfeu2hWNT2FXRAfSa9QIIDvUy15FuMhRZVTYm7vHqfyY3tguyzpFVTQpVBhaLWp5qYWuZpvuGe
YWPI0DrEfkO0llHXr6d8vrGcZSSz7PGxnMVYfUO2SyMQNH7VpnAw5gMgQFQTj2FsY1yXob46fmZ6
5MFXz0omuwXe2JpE070NQ0nWRq+6dm6eRM9giPXDGK4TUMVcwjPU4crRlj83lHK2QqTNhTX/MMKI
ikXina3vlEy7gZFe1DmNm/giSe/7KAnp9/6FIR5MSHieVWsZb+kBz378RWT5iTkeTFiB8LkH15H+
wtDq4810+AAo64H+92WHAeMJQFjytmzTGgyEL53GvpAKgBFNgpovPMkDzkvYl1qCSEz3T9J1Z6pP
bAZe0FZOy+KWteXwNdCPxxFBblRrhCS0J/y9KtmcHbmCSk1V94MsxUi9j4g8h1CZpvdvGmQdviOE
kLBn+gzKLZ6Gt31d6ZwNv8zN0nDw61FMEKVn4ptEl/i8XfKSk11tKiKviDSfb+2bEhc7XG8T6zib
HvDv0PDMlAA2/rfimMUvcAHBAvHHEM4QyfyYuvprX7ZKrr7DarBuWIazfImxal1Pbk0FHgMh/tW8
JYuRjEre0Gi6Kdcr3cFYxI71snDt0q08sEEjKFglPJrjmgwmE6YBFV6bLs1ChSeUDWMsblA0o/iU
gC2+cTcwZJw1BNKKPygvqtkA47zm79MQX9dcCjclQbiiN9j3lK9UXwB/0GnT11Q7xJxpboFuxn2t
BNnuE57oklxy7932orjR+6srP0khqCYLhwPfHnLC7YCxAQ3gAz5tqvaNJhW+kqz8kS4OP1moEG10
z3mSttEIU9RtvlGlds7RYd5EBRPn523dZU9GqAZVgN5YksYY8So8P4IR1l7piryBeIp5oeVLUUbV
/Iej08bkDNObZZw6p8chI8AbPnlSeAgaHjkWbobNxrf3jN/XrdlZKaEuErTshwRYRyJo6EgpbfEr
D2jc6XiYD9DXtqg14N+MZOcQKotIiywyF4ppYImlsfBuoFETUyQMZYUqluPC3Ttp0GXBZACCcaEH
0hBOhOMFUg9FRZyV5C5laxqewHt+yYDqEN0RZt1Epr+sjlS9azUU/lUvURLaR1D9Cf9eHhMHw5t/
pD1JZFFtIVWIW/ij5vVaM8k1Bi/KRhjnl7qWe9aGBBtigggFz4C8kG+0paqN2eFSHArME5Y8Ta8p
EQb1diXkd4aaZ9xbhfqo2wBPzHP05BiOkRH3v7bodf+7ouyHzaZ7QPMlPABzkvUY1CTa/ZsTmRJv
RKLw2lMxVJxiErbngRFp/gN4u0q/2WLIajT/qDuvn29UE+iEOXD3flvxjE4CZPDjgp8gxupUKPSE
XrPjCQaPJw75ARk/YvP97Caiwk8hciDDPcB7kFtRaV+wyQPfkUwpJWuSGuUohjefqfgpuDWxNWOn
7m5iW3gxVKidrCVODE+xZeGqrRBCoq+JRdeuv+l8p8u8xLC0ExKRa8fo3C3FySWOzzMJzPSlUxaQ
o3MYlDqCMwIkiMZi07IIW48Xn+TgDi+Z3sLVSdxxuDajAlNRwolB1pdHDOJYQo8oOwh4kuH5S04A
o+DerESNWOA/1jIctuPiPhvNkLeW8eJlcvI/iJFdiTJVEU6UN7h5tz+8c2IN/FrIAF7+qCHC4mI2
O9H4qqE1P7h0Bi7pqEavxBn1LoUY08WwJAPgPH6ABy0pr+7EZVwr88BwzHhks/0Tpm8IymAEMJBt
jmfg93/pzzqjgHDlcKLWK1Yg5v6vyFxdJ3sey1txG7xvcbCdJpT/OrZ8q9r1G5mK/YVWmC3owCpu
h6YE/z34QUFZB+1pmUVhMp4WIxShwjnugpENRsV+3wW8uwH3XDrsARwX9IeniupW7DQ0H4NMT4q8
h8gIgpOj6n1boYuR/1C7aoq0DsodBL9z4TV4zeixnR2TQAU6Yy6qwdUa4V2BBxZ5mD2uJIj7I9K8
6Qckus0b6IG9V9Rnub+9WJyhNKzbRLl23X6J0oMJC/PX4MqW5mIlEkduC8SJWLn0Qf51KDM3nNNp
cvMIyk8JffJRGJ4yz+868EGS840cy00l2MDIdpAEUvgtx/7joB8H0ynUx8CyQaCHUkq+QmxICibl
676nPmhFLbJsIPrOdtIIhFOimLcFTEEjE7uuaGLCwiKiyIRw1O4eNFvfICWdGLWkJI1k7/F/Wi0j
dxoCWneesB3WPoXDt1YIipBj5liF6sRY/qOyx4gFLGFHmdcbd9ao2/zcudVmCeGeNICuWxAYQF4o
ZfX6xeRC2Ud4u5fptPbGjxus1AbDd4mpJ0igqpa1ywTN/Nx3BCQzD/Q49jXa8B+Ey1LoG0OlQuFh
GSFVf021IQheDNZ9vdgHunbbtEtTIhb3gctdLmo3sj/V7fUZgTUzMrFt+ZpGYA1y5Rf03e1behmo
kFT+AXERB9B4WlgVvkxieDPiGb9yXolAN3aNBhGQyIZaKX3VOiDmO+aeIuCqtOoSoYP6WU+VPQFD
ZUxPObplOtyVLynFBYfr0ZZIU57baV27zhtsT4c32OGZWOOacx2KaTFQFpUeEMc3yvdHYGY9ngMk
toK5QyCr7JgUDHvGxQTzHpJsgbLusV3r3aApR/88Ypw0bKvFFJGerwtDssFacsiz0Kp7rQB2++cb
0IHOs34SBynhWE0eEzm9KHEjWzci2HAHKiZeftM8cqwmYqjcyNpex68JJ+2/n0LJd4Q1jNnIAbp+
qo/Ff6ZlnldV4w0JrtjwDmVBkw68jBMjNGozc0yrywYAXUyJethFrtN90LlTlHwL0FM/O8rpW7Q+
skel06eGrgoHROdbPrJmfwbXkHVCXtMIZgrzISyTm7pU5IIegEd7hOx3JMGfuhe0vCfiRlHI4202
UhjfY4VcEEQk3npOSU43R9HAh6wp9CYtGRBKXj68P3LL1IzILqBoRjSOoCHIs6jisi9vYtE5VPcG
K/x+jwFMEJylJuoG7tzFtqqxoz3vptsUugd11Nz/digrHrAVSuT7v8cxB8RokxizJB6F8rE5/XcN
BW7HgJnLlIHS8QNMD8KlOq6Bnm+S1fhPaiNRKZSpN76WEit28W/6PJsFaB7IennYwI2jvP3Wp1dd
+pfKgrJWk8iP+qQxsoDLkzUgRKygcg3no76kMt2SGWbSrn0dnZ22whHNWqz9/Gjz0W14xJj7laWP
ablpPpXYalRYOpRNAzRwg0CJ10HX7oJ6H4OjELIgVsdfSLYsen1XzkfmJm/gCZBMOy2b+CDVast0
paXd32Vwgylo2+qULlFFxPkS6CpDDNxQoL8ss+ECI8o542UkXdEIX47wbmM0TrjFZpjuK2Bjom7W
22D7ZweQMv/Aw7H3WjnUEO6ylG84Z7o5bzZstgred4UykCnSUkjwf3ho+XL9BHlK5U9IVE/RgvTM
4GafX63QEOTYVrHNZ6MrfUZ9ykM7QQe8rSQvdfJmTEu6w1KtRDo1nJSxXeI9nZy1DnQGVZ9uJ9OC
pm26YH3aM3pmLTrX0JAXrp5tqOB4BQLFtdR9YbA2wQGWKzZ7CbBL4HXX70a1CbSMaUmykVlmMdjQ
OggSNmuDJhWPyRdSE/jdggMkVMzz9CQL3/RkAXIy7U6svqMxuGNEr//yjMZdziswBj2BRcJmJaYL
nRecQMjTDd+ZWFShThSMmWTzV51/cWXfiLK6L0RZHWtuEC9Z+rtIsufjqFyz4oh/KJgs8Tyn8H8U
amec1t6GpFydDcYUyxrzo5UCL/nN4QpYrI+54djNkdLXJWW3wcKHBnXH9IIJYZ4MCqcsVjze/hYM
ZdgX8Arlc1oabFZgVokRcwZ48qkgyZxj0NNJT1P5l5SRcFDLwM04o4CjxmoB3cjBFNTcB2GPZ8KY
qZvC2VD0/OBto4WQHhE8LW+ceYDVLANuyrzAOSqkH6imfqytCqGD/qZAP5hmJ6SHzgCcfnQ7asbH
H+zt3SVXkdG26qiJ6MZUKH4zQZ2oRbOxNkZDCJRs6c9HLbRSoVMhwGt9WdgpQFVzEMR4iG6I3xMr
/OcVzKPtlGkIjD7YzG5uEK5e5zXrxhIQu0nlnT7rCBeFAvRxaQvvKbG9S0/Gr3Pp0GTozfL2MwjX
hySUqVAQfU5VAhDqOPFRURhLKoQXiGckUSQu0+jXG9DHeBqn47vzmO/QIjJG0P3dZUBpxU6dnRmm
tw7Ue36Y25WZx1dLHJ16zT86ji5YoaL7cNGfgmlto0iE5sBUgfkzwq4LYkBj0LA3lKXwMOTXFgM0
LG4y/26iWYzWy0w62A6IN0RkLqzvqYBWHFIs40vq0i9CvF421Q0G9cwFa98anUAtJI9RwB9a4UxP
HfkmyvZexxA1sAfO6MIVQ9E7a2ZOC1RkFME0jYl3TNaNAJ55/uT6GMCehcjfBYDUwDNmHc4CfhoO
dwnKMevFzeo/MlG+RXJO7/WKIfS+cxurUjCPoq7mOF3JxCCIrD0j4BtjuPKdcuLKcTNVapCZKZ0D
3X2bPieAvikTMGULmTj+ctg7aibArZFdoyYDzifZHu9qdjb45Etf8qwadF0VRSgk90HbdFjYaDR4
V8/Y94waCVO6BRXGOA1ACtUNyHgNs0ffQbhvL/nSAPLEVd7XCtDkJ1KUice0UWWzIqy/8rXLLsou
fhhjPnMYJQMZlhRCwxv1o9ktVXWPebohYsxsruOAPW7lMPwrLJsEbZnd0b2X32nnxgP1dGHpu3I9
ud5sAUEpJUgIuegTSL2/M+D/DmUdJUoXlU6EaESDDZU3Wgo8MRGS20Ze0UDGhPhsB/UHqlaK4OA1
5mnsnMHpq74+BcJyTjWg7x0HwVuwsruDEFW7ivlWjXfgVsd4gAMNnJu6l9MYAGf3hQmcVeAGlqmT
QpO6ceZjELjTldgC1CFHB86ghbs0jKaHfQAOgurtgPRLbkSTiC37NN2UoXX1pIV4eBXwXS75EN1A
lEnDLVZ2xKYHb1siby2K5JkkgtoqrriqhVIRFHKshbKwnzWaipV9dc1PhgINUiGe/c3aSESb0S/C
MBkW2K+HHwYTK+zzjk1q88XxixO2ZvZfDVOe8ZAyh3OHWY1e56cUPbdDV/+C7DKFCgz3MNow2iWr
LcrQuds/ReTN1z7gFdptbEBhYde8L4lVUs9PJ20aJ68zLPqaM8nORRQg9idJGW4uQ8/hofy3xKD6
sf5NR8A3ggF6WnVbmpJ40kfeU2Y7HxWrBXsZn86b8lxHA0Asg/cPqMLY9TGcTPFtOfOJEepEncjf
SAiqL6x2Sd7tU1glwtKQojSzisz5A8+2toQuQoJm3rs1Yr4mepNGAce3/IMaenHR2ajG6h3Iie9H
XcSch7d1Un/Jhe7siP87Bru6650GfK5y0xZpf2Z76JVFVfFU/YCw2CQCHj8eOaJ3GArrM3DHWBru
KVNCjx8wgiBzBoZkcegP3CTnNUN/0pooEaTTQQcXiKdXNhJeBX5FgyW64iRVhC4sydrUHOc4o+sB
0iRwLnUdntlh6FJRcSDQyEszvVog8uRWGbHB5CSfGJaZZrUV9dL8IFSyA4rfHL/eLH8IAcO6JL3W
4Jeq7AnSRwhz19juyGfjhxuQ9BH5ByQlqQR/OH11vMUb90tP0Kssdv3+b2lw8X0Ym88sObnsmOdu
ZyYmbE6jD6+VrXj1VcOCkiKH/TyHAujCdlflxTU9cnQqvuRM3D3eoJmV8TfFDXh1PIrg8YsoAomV
s9kpQ/VeIyWCsD3zRuK7G4CFfenFFOeslOaR9cOlu5QwgdvXeasjEnwoxvoFD0TtPJtWJdmk8mFJ
oqr8O3AcE/7IbJflvMqDMwEbI+8Jt+YIk135il5lyQee9PXth+JxB5EOrB7ioljTyYxlDT1sURCn
T/AR+UcbBPsRazbAf13K60woB2/DXcHwOB0gR6Q7ob+kVzSkXelQUZje4L3exPCgJEvVXpy0gw5z
lJEaRLtJ/7Cy3LK7smzl10i4Mb70LrYwg4hgsR6w/Zrv1n9HTgefkIQQYCSk84lrRK9li6YoSxqg
6S6u89Opaevi5P2CT1JsQcGaGKtJPpPGszppd6LrwjkORLUaIqA8USLIrcBap3dmzKJWTbomRlB1
n3njC4ckiIcFlmEBT4TPE2f2tVprGL8N9tzEseq3MmjtMCu7Lc8tg1GjxG9Ouexzq4JcL0uSamEf
awlmxirjAEFMQ88EJ3xkHVpEZixxCqltCFs0Mfwxp699rcTmX3TGIxjvEejlngTI1RST+wivhleU
wnCVhgSgT72ryuuFFho+9TOZwTtKCGg2ZHc8tuonX0kjI7ZNzNIhcNRUJ3x1zaHUm6E5jhcahwDN
mKCSS7xttMtX/v9snISQDVnkKvA9ASzQVyOMqlLqn3brVArDKKww3RmfDPEzWpF62fti+RBTzQ80
WjBDP1c2RlU7OxGtantOaq02EcQU83jReasFTZYLkcCcl9ue9dtjBzQn6ofpuASt2XOzkIKPGj1Y
+NR5LZBW3Kl+cTELSu3adNEUdGxg/bqGx6knPE0uPGURICpi+TBTmcyRHzowS4KtThLtA8FiXmg7
QU7n0hCisi4G/UUZVF965HKa+JZgoFeJasso58Naf6ySsM2i6d6zAXEEBzpu7bYNOvOtwdbhJpKE
65kAFMC3/gXL+5eJm6qsCS1HCijnOdIPSUak+vYPgp0hUKLO+zWzXBDsN5wpxBieRBg3XKU7i4Yo
nrVnJi5ZyZIaksueMOdcMk1J1TviQAgZ2fyLvdY8SlKXb8qL0rlFS42tdAUPhQqugBTrCaId7hCH
iHq/fWKpCxtxk8MZFEIReaHya/xEnNxCw42j0YMn7xP1iaSYeKzDxSrg8PkpFkWs/c9a+cebkrYA
VJRqcr6Qv3YFzwKRvg9x3SyPydEvVx25CkHwa6W9OPePkT/QW1FhJnXyNlfDvXXchwZsBSPsS6rY
tCvcYLe9v5GpkXXeeYWwVYmI+Pyl5i/D/KDVKprKCF379Rb/DuKSNpMMusNJGyhVUogNYoBsMXXO
J+1bOLY+Gf64uSD63C0KviVTsrvXGYmGIs9m7NcL9z94xG4D6iaVdfw8KxE2kZ2i63HztZAqU5N+
4UY8/Ld1QtzP9w74V4okI/b2M2iG0HI9+GfDZsi1w5fW/4zjrISBMqx7yrU/zFDMkzLZ0e/l8bwD
FWybsKjpsQ++m7e5Ng6EgMI/8Owgl5Ka4/wuSgeECL88YaU7tm4m/QaHEOfiV5l5ijDXO/wKQrfv
8a7WueoSJt6AeJv3CntN7Ta1iu/s37HsvtBJgrkMy+aTi0YrI3IF6lywRHm3na4qWdNwtOwokynV
9afWuXL1DTFk64ecC3M6aVO+q5KnWw8PAjNeV5ezeav0Kx/9HuIb2iadgp1047UqmIJpai4qUaIV
T60vKpydjRQR6et0H/F5iUHWyHv8hNnlhwoaBPYE9L9mFxHakfR1BDkbzQkDX7waq1AdaBShU/d7
LQ9pNo0r39hjITdgMYJp0gvPXDLprIldCcVBYbHJMCOKoQ3G5V11p73eajc729p8tO/HHui21Sli
7rVQ5F0+oGvdvs4iUCrBC9yae6sSJboiphwtTc2hVTaBsmGVP/J8HUStGBdnfaNlqXfzVh7Aqswo
4Ehxie9qjWrUvfvkqAHRK3nq7TzaoCUSkI075iEc/VraR+TXFZ9m+HrkOD4ezue4n90tfx9MmczU
u44hPfkMdP9ESLV7lNXSsus+WcRmXuUv88FTGqdoJcj8QTcI7kXtLj+vxZnOlZcFergVNZqEbngx
uPMTf3EOzLU2Vr9FDTK3I9Xlh96uxT+c7Jn8zErqpRz4+SxOjkczAueBu4ohN1u6jiwQcvOM634Y
md304Ws41XYRhfLFY1PD9mdOiofqtHL6lXxDWdvJeZRy85+dsQu/vdLJjpV+4dD4jE85zaFBfJ5j
5tkhS9or54Rps3MqIS6/uHkvu5jLz5jsXknn0rYvS2jQa2JS7SkPRclJYv4Y2WMcyT1hAw993vlR
mrv4jxpcDpwxs5pHeX50oho+Iik0lAEix+2GI64J0pA80kpjS/TLbyUpQ+wwfW+Lkko9QkxtWmAO
xzlw7uUSMHtEZLNYKgDdR3DplK3N70OQb05Ov0AsNsrgPN2gLP+1zoRIWCx6SqQqoz4ePhF0JMqs
xJisLWbQEwD4T5+YMDakLmBzcdHViDeMrRmaRiplgx3HUATPzWzmSzrnr2ee8QBXeWZ86d08Up6h
2oelA6wHpQgR5kChPee6LkHl4MVu8LeBEvwaxp3m0PT9fIqG8DHC9mO/DxIPmQ301g8EipvxXOCA
rFJ2mPgR5z/OBXd8BSjvtFWMLYLiRJNI8x55GWkNF3b5+tQ2B5HeODs+t1sWeK9cRxNvcirAEP14
ymudhbxFOeS0Mg0KSVhxA76yjdxNV/beAiIw6C9jZv8T1eJfilq3nVb2Ebgs5DtJgVW6e/1RaAcN
ChCNIl2jHBciXfWBxycu9XMbbdYfOj2PhqjIaxeDeu5yhZk/gd51oh1VzhPDtyzGvm8uu3uFEAwE
Du/RuookrsZBwM0bRNhBhRIELkm5VtbW9tJfXoD0A4qiRtwHN80lPM1wCwVjQNwEf0K8cPzVNGOZ
dPu1ldmtjR48vhpF9s57aVvnX7e3HHQr97UlBtO/CZa8cC+JyDPzzhd1YhRwuG4KX8o6Wv94kFW6
Q+slzSM3QuRKbGEFJpJXnt+KSAn20G83dWYIeMZvEhqPE/ROyCRq3ZLtUhXjN2KH+4wq4JcIXE0t
E7ttZB1NCeLVaqE6aEHn0KPufRlhFDF25GEokc/qNCAOCs0x8anU4ice9dlPILopX2qQBEGpRQlB
o82GyOMNhq5SH0q7NKQz6lnVrUS6Zy8r87amewfG9CL0ejfeIMTmuCyMjATZQ621wTWhebupQ0wd
YLITIETDwm+hVE48wfnrtPXUYGOd1vjTCgIzYZiKsDBS7O8w971pcZsPoSOf0oXcLHcYmoRIu2Ew
RlAdykzzVh2UneTtYATum2Qt7zbrBeQXp9eiL6yg7TZG1bF7POX87FnuHCXHq7DNOuMUpMsoPNQ1
Ly1nYm5gB2Hx+lnAOrAbexUXRwXpPKzA9JqwB7yxfaK+JD+XCM6BZrC/e+p44/CcBkM9kRftBk0T
3o5rI/JXc3Q13rgewAwksP+FBJFvB24YDdg5lkrrqfyHTlwE4HoGUcNIxacjapvxG50uP7fOMBMI
sn75Vuo7wW/MTKIZdwVsUNKPfrcz5IJZtU63ayFdl0sgBQ/JNuFsjgU6t3irndhX5bdq6e3vxUHC
QvEv7ul4tEytJAz9bLZ3AEV/bTR+qSKyumvs8XYbklysOLKfzOu/WLHwVKnZbm/LI+Ta+Z1rH6d0
8PCaYpbEh9OkcSN3BgZYsm7ZavOLjKgr9gCiz6jh2ZZsPdr68CPGGTXNe7rFr7MIvyjBnBfkwQGl
m0ekncwkj5dgGUQhv2WiOF9RB99McHcmqsIv4AiZBKcUxRm9D9lI0EbvHcEHx9DlgxqumBvKhsNt
W+IcrsYKy8/809tbGMLZuodsDtE2YGSyyC7FRPkMjvcGtGZXpgjliSN1BNMxAii2nQkSipvGkad+
Z4tzdRuQOd8DSa3/2vgBV+IMY3X5UC+Om07h/AmS+K3NUIyZ1p3DQwNdAiRfHxeWzw8rG9Nn3cDA
UObc5p2yk/RTixhUxGlHgz0pv4oHIfF/ucI05Qaj03Da39bv1Eigj8fTwyQ2upmUb/oqJdfT8zuX
Wj9NMuk3/d18FU0wIzwDlr/x5hdJG1Dp5trXPB+CSD+ZdvLrKLYmLUhS0YHBpcHEO54HGsF4UiBL
KNh1eBX1GiMW1AokQpXtqP8/4oOtlPldL5O/FwZAQWkkYd1/eNKfNZsBlvwnLLyRi5c50bP/vQqQ
d/zu9U+x8q+g8GaFmciV/ADKXqHT1+aRBMlcgKmUfcSrHJVHcAIvCnJ25Uijb0w86Gb4oW9qDjIG
9m2xRLHW9dINuTSpSZeD0hAq2ZhbJozZpzAaVqFnwpC7tm1ze8utojOm11VeLs67ZAirwKGM2Xcv
nlovn4iUrxxPTBLt5zC+2QZ5tNBp6nSguFhDcNR8jBPhrbEdvhBUXNTk5wbRhu7E0M5h1UZUtJaP
UxH0ZnngiRkV3ff64Pz6WbP4remC4JUPfGC48u1B37px+tdzZaNhoc/G6i1trEUUhJX3CAoyxVLR
WptKymnShDe/i7mo4ft+pahKUibjf5Ns1umE3rSnmycWpbnwyRE0sKro0rA3/P4wI9qHlKymiTP9
e7b8s45bbcUI2vxXVwjt4t73ruHWVwo0aAdb05vw/yxoYf6aIVHuWMkwmt0H978aZWApGaXF2Ce+
WrQzK2DgFh/JvuHZi8aqczv05LION1rN6Ok+XN4BbXSRqRoJrbWas5H34AFTGSUXrl4DhCw4JTDx
g5ZINiMnF1Rb7UBdnNL4RFT1uf53zS1uD7PziIQTs6B+GxI/KILp8WtWM0a9Y1mrttA8D2f31eRM
i2UPkS20X5L6QGXLbcFGOmY7lS1K6nFxmTLbZnqecw7RAqsl9UjBbJy0+VvEx/8n/L4MHyKlzLLc
h2i9JBvXDq03/Mnx11GtySYyba51kKVWLGZbVJtQhptDxxS9XF7YbgJUCMLgCcOTBCy5NyQV6EdH
Kjve7yonOXC3P9FqNgUbaVRxjBdTDce36CGO+epxrPOtg580Rv1x4pVU2JkKIq7WVTY8vK5749w2
jggoaCdfweZh8NNVx4MFZ7QMbOwbbMoeklpnNJOTSh1e/ja32/B+DRMqqR6RQKBZe/sVdaaAv25+
ie3XhJm/tqcebsJi9NP9Bl6k2lpKqs06UJwt4pzY1KJ7y2Ho3kVJp8YOBTIatdhyjiJjZ/3UE/7i
WZEFyMsYtYXkE0kzVrtbjE1vVEOdMjoOzPvzJECy8v9OBhdpaIh+0v2IVhc7yoQuRjGX9o95sTto
5Phh+I+KV4zsz/FJ727j4WVe9czxefA8Y6R7PA7SxUuj1Hnvcsf8O+MFDnT42+QUVPkES+B4l5cS
8Vmcm+DDTUMokCujfIU3bjwRBjbK6wZX76OnMxCmDiLVWB/7YsgWHfL5c96H+ixB0yhiT34/bdnp
2tVNS8Pi11in2EDrdsXvXYL9IGxe5ueqinHdckZL3+ZARNIYK+YmZ4T4+/PGwFy0I05K11zZUJtF
NWwk81dEAY4OpvWmFvqw8NtPAs3LDatQDGxYUZs3slJFHT8VvBGFoe29txoKcunM0Byvfw+O0Kd8
UUbAa3FIo7rgjx/BYzabSG5UWrvNEYuoS70yJTQIv8PZigmQzeOaH8DHRl9znMqOS39PHzvuctRD
zfIkuCgkCbthL9f8ColwJ9swpS8dQXfWvHnq513tN8V41+oNItElS8IUbyJS51lDzym8V/swMvkz
Lnpx/YNDRMgQMWqOdAfVyJcnmQ0qlGF84h4mua4f1I9qhHVugJpAmAVphLwsQpjYfE8FvNlck+4z
wndVk1uT6rnGh6b0NpRvcEiAYL54LS569vrBYhpqbIMb/VYNaPyqg6HYilwLutJYH5kRZ9oJ6aSO
uSBZ2UYeowTxy6Ww/j+wyAk+r4sPI4oIiT9e6nWflVefODnKpJ9wQIcXBjFgYZ3s2jmwLyUVHFI=
`pragma protect end_protected

