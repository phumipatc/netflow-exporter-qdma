`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kaeveMkLJiHZ/QcQT39JKYUHZP8mfSD29mL4L8pX+foKJA75zr67cYSduZxkJq+3q6b4KgX4NzVf
CG4epKG4o3vYW5KbBCzlqFqns4CN3sIMfnV4p6nDU61oKBsiI5YO8RjhuuYwnkOJeKZGT5vnW2HA
kDxDu5sHIYE1ZQ6rUpv9dC+sSrsNsBbKH00YEz2aIMgUgRogaRjC+odWOcWAl3gj3Rc4sVj2qDWR
F4m/QRAqT7zX+nfDbY5j54yBo1pWNhawu7zTF1QMw6H4Y1QM2K7Z7ZCnWxfLamxiEze9YUIV2tC3
8md0rEcFBz+MXl4/mnQ7qoIMfhs1JcgB3izwtA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
i35Dy8WpZ7BRYCNNSNiYDgUTCkdWHvwrUnjCfarz61dZdvpmNCiFnjgadqnaMka4MeJjcnNPt5gI
h6jtqA7gFTfk3rM4ZIKMsgMcSeKrSt5637PgK3txOlam5TMZUEX1PySh8hhR2bUcALF8a2R0Vb9/
hGOYBwY/+a8h8jEHc2ReVyEqe+YOBWH7jBXoVzd4HkdRz+JyDYQJp61FyzTrPqWjwZTxhyasd9xT
KKCc6TIgHk3WyT9IOmTWEWGK+FCSLnigykOxsT3Gc/nw1pH0PIp3YwDxm+6BKrfoLMxK9RpXA7dm
mUNpoMVGWTlHenKRGWqaaV5mYno6uAr8zOJAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
PmyO9LLJySrU97WO4fiPhrdJXMexCU41ljT41ikbuYMnvIJkyyvZz0+kYbfxHZtN2AFUZBslU1Q2
9O5llwB1/Q==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
IZqrziCq2hxsUgjbX4l9gS/ZAfMPw9h0a0IPQmckjfE6IGBOyU8tn8KBCtNg38iHyQDHVNJsTB/5
dOMNcYv8f0tutpGZteXfBxNzPArUbk3qVDCMqnfnJfrdNrBwZV0PE6YHFO+q+1oVvQEU4+o8MrEh
ObKvQQ/mrFfy/jSi2f8hVYcR3px1ogzmhHsCrfUk07rHVYMFnbP28MZjDHORuSmhQm+fgMmQypJH
odO0knXXzlYZ7em2I2AO4jApEvjrRHgR+X7TNBDyVwkUFze5HRgTu7okRs3GMNej7xsmZT044PSJ
W1PxnVzXKd36Ek7DMpiE+njhjdQNYzUa/rhFBg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gD1lWt9Eb8qN4f+FVcSWIxXA1fEjxhGxNFyg4/lGHkTocObM4HAbCqRCfE8W3HfHiorkre/0wHdm
lKSLCAx2kVlIR4z7AnQ7bjBwPOQ4tR0z65sueXTmFD26AteWbF8dNRNZZwboQ/hkjdNEtlacsS/w
PF2tgIMwKkkhJ9zhuP22kqwnPPg0m/mTdC+IU6YChKJjlQfpI2L+D8N/5XpEmuAI7/T4HL/SPznR
1ZMS7BjT/dp8ReWDmlP4g6ISq5reQAJYBaT8Z5DoQ6TWwf7KNGrgDrsi5h/+mewd7NU0jmEQozcd
28p5zh9MBvna7/Xl17w0eX5xEwmqV4knzkpIpw==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
OJlw/AT4Le4E+0Smg2g1oCENCcvx/W9jBPjuKOy5XuR8LQEghNMZV1WmpmhuU2cDN7eTQatb5XIW
0eRkcIeBp5uBJ6EAl+B3E+IEq2mF7r8Q+m1eQPbhc9xr3EaQmC6zCwIBQ91yu6T0jyZls6mY09MU
31FRUUePmuEytOIkL9s=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Z0XxwfzvMXyy1C72JWwKP5h4zFPkBJ7KXjoEQXPNvWZ/SCeClA+59s/V2wHQr307kjK1SgCkHGar
zmeBE1ZOYnpSVnvXLLrSUYGYNkUoPZcclreyXaMoQKDMFgSBaRkd8wJ7/Rh0OMBB5Lj9tw0SjNmx
qD9Hvxz1cosLcJxJcFwF0NPDIBVsOP3BHcl8Pv68PAUz98J+hID8XZHpIO7Vzn/73iuEexMjHO2X
QKTbk/VzgofKXTc6bFxzlUXBKqqrwyfNEKAaAi8H4UhNwN28yh/86bPswsxIIcitGVWlZz6QKHOw
YunDx4KJHpJ7QQf66/kE1+IH82jpaiaCGfzfEQ==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZVlkl3sgb7bW+ZAOrh8SNEqTkf+PoFJDO+LgYWOTDqwR2GXANFNq8D5FOynubqaaY1kp8QJtV8sL
r/4E8m9zWBwy13JlzFLXJOENw+9xR72+RnQ0Har6q+zjaiEFXIHlJcns4jl6MFSJeo/r6f1eNT8x
hOwolV1jV5gBqiDoHNhd3iwq6/wDW/htNdaR6Fe/Gs5lfWMl0w/sdRAE2J3Dwla/DPQoAhSgtb6P
/aYpXqrOTRK0so1x00RT9KC0WXBO9xiGmxPdPlUUU8m7kcbMKIJiNa8IrM71DOKfFcrBkpeq0k06
AR4+1PL/ApvNheshz36qszkkWjQGpUis0gw3/w==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
u2gnOuY92ta3juKiGgx56l2nVsDfJiWI8u+gzlWXiz2oxFU7UXoChviO+y9voj7UsdI5FxlXy7O1
Bawm/PN7hp38EOVcGHWoYSFNf//f164+YIEIXIP6e3p2z+9OJO+5kxjxxv8jZcqqN+3/0ACe8Tab
WgjwpSlrn0RKWVpLD0o=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RmX0VPNJPfZ18qXeRQ6SUG9OXVvoSC8IJmqCOyT6JA2OkzFFevDAmULxkXyR8yyl3tvEeeoSo+dP
+TVxmcstaBsiAGHjCjfEwttA4iQ9SecDEtgawZJ5pC76Wl1D9gTkByco+L5lTyEpBD7m1rqQhQ1x
JrkMTZiFyvDscBJ9MBIrMz45c/dSZwqIx1oUXKQPTvtBKlU1jc8UqI1+koNy64YByaWVCWNkrGVS
VAIY4z6mdpFScyFxuF+Qp/0KbivL8tRbGPTFrqMcqubUAJN4LR72LA9BDdtBytkD+uRyOl/MFKTm
XYYfn0Joc/ArluIIZbqbZocNagJXjL0iBICbCg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15648)
`pragma protect data_block
yvhQdJYcRCngZ0FBDXG6J/6Nnl8BrPMp2IMRzK2NXQFaj2+EM/60LUhr0MquNSc3Qs//SPX43yp4
4uKua0jYvLdW/Zv0CcYgsh9UyCxUg3zg/kcyZxqjeBzJdJMcqogsgqdgdAn19BKSI9xZaWpYwcjs
d1dGRVwS7KjPCktZxer+ngSUik2cbFF3orBh7dr0109fvBV0ZbZlfrt7gGSA7szexGnOA8daV/7M
DmjDJeDNdKQpiMHaSnOF/jZ9n+GnKF91jJlhrMH8HN05OcCHHakl2aREsz7IFJbv5LRlpWJ3vRDQ
CD3EJrfeYnjIUb2UbQ0BRYSPRDN3x+g/M6vr8k590RvVPfuoGNCWPF+z9PYaXZH03MQEJPNZ0Fxd
5oICZVlnNZezMVop/uusHqbq3S4wiEgCEpEiwfDjq7fgkMzw3lMA6dLj1J7km6WzZkXayaCf3Wqi
BEelj99+iOjsgfqw2sd3xQjUw/GYyRgAtnJ0L/n0XsovvyYopQpXdiPjepIr+bo+k+q+NQ0N0t8W
ku2KH+XRPIkFiVCtbzigUPRx80lNzlqTw2jCONuncS88Gj8e4VI7pcMac6XWK3f7lIunT5AeMKTn
9+6HbJwve69FH7HwK5/kS/s80tq2ixhjpku/ZESHOHkowQAfMWBA5WNozVv2UaVVeut1iGZXTQ42
iB/6dbPrK2uEIlfOMR/IzgtjlVYm7AyNSPSOzNLT5gwZAKIUNoXxOUUxlMu3W53rv2Vu0npunN2O
DdYc1726xIZ/qBTzVmouiLD217r7x48/uV9LR3uJiKnNqM70RmfHdUlN93vJLCrlujXB5IThTDOx
zjuB0SBqzIzdnYKZfTxXvyQLoMX0C3VO3HfIMwMpewSKpfKkKSZ4LFK1CIdmzs//zu9ypOqDvqk0
9xY9TlEGLG8033lcn73pbsH1Z9pbYpj4IPYgkJ4oC7cbI7uOnUIx7dDM9CpSeg5OdZLcvz39W/R/
1ySG9j41Rk/sKDivhSEJGxCSgYADXSUzJh9DGAvWKtORTuu8AJ8K06WAM8CyEW8IywiitO4fSeXv
i8E2RsUwaNcxBDfxQWG3QTnk+mrAjvK+zleV6cR9vCwNXrBdZh9CvfW4YelRCYlECiIXKLnugdQx
FOinsc2q0BE+JwzT6KMaIFQbopA8DSiXCwULAxyP+aJOmWb2ijbRgFs314TGisTyfOheD6Wq1vA7
B3STzgMxS2ICqod7AgzBxWZqvjWvZbBoHCvdnOFDauoG8REnDBEXaURTy5dhiAIdcxKzihjgAj93
P8dg/1re6z+SY0l+nOiSoL8uAnKxQXFZgI3AQp+67+3+QDb4cZtst4BdB04rESLv0vIMttJsGEn0
esVNoMeEGb4+B1RgCTCWoyYO3G8oXTyrVQJYzGDuOjmXH4zjSs3CC1mbYlvnYfkASxMMVpRt1ZmM
g1IcGYL3qLrgIQhLNUbebQO7U7+cJvxKLWMg7bvEXHhexeuGjDc/gqFYYrqRSRY/YkQgmGS8z23m
onM6PLVTH/DZlO5v5RouXv25vJKE5OfjR2s8a8wXX5jEhUHfACTCjAN8AbXDSgxVZXHT3b69zRw/
3KfhNlo8FXRPstBsmawrZ0ZLIorW0C+J2XfXSL0Z17RJ1l4nAlECkt9+Zhs8zIxBYya0cJKREEiP
mQnYVG/IWt/DpxYhlDJwc8FhTe9hVt+yyH6oLzrBnukcJhpTLCJbR4JevU0pmxl7hok/YP74QX8d
nKelmgabntaIqFDH2uvSCPwRL3uapq3n0rWP4TR6OLvKg2TPdNjo84YB3I+wSre4bG6lA8WWXvZR
huVV2J1CjjvApfBLLRinnDfU9+WAxYsmkfQdjkoPG1/1EC6mjRapWskhhhQ522ucZrk8SlmDPNut
U1N44bvxux/mJ/o117r6jDXZywslI+2mEJHnwQ9mWm2rgUIPP+LqpVqYJml4o3LoVdwJXad+TRCJ
v6HWu+1oYVLNj3vj24pMT5HWfBfakbGphezoNW7Vt0zz7Olh9pQCUfvtrqxUX1Wf+QEs3YqqJWvj
e4QQY38TFPezj5C0J/jucoSctN3gfUmYZO0VXjTOf1I52NVIpiBirMCt4y9yLSdqpLvl5d2wHlVK
ILjAeRBs0NmUN4g2JJBeOhLNncgpIxjD/R8hCC/H6a0UvMyTKQW+uG6p0++ZGBoCrwggcRT9HHCa
X7zbXO3WpnrnnhK6EVsAneIMR0c6MeYhw7avtdarD7QTSFAbCpvm5phGexAfo9lfBPwqLbLAAQVv
fyrNXieOpA7o76OBHooY6CEQyMBi9/O1yfkXi9elZ2u1m1Db8w13PDnBZd+j4Wv03SjMe0L3gXXm
zowWZsLzRjghE1BRHcEfjf50tW3dmPPRw6hXxjRxhIittbowIwzERizDxAi8X4zYk7LHcx3shGJ8
Ek0RCJiAZOeZ2P022vSLQ8/6B4mMw010IXoNMhCj0pQUjSwpVgwR5FfoMLdY8GUZLEE9yAvsMXi9
GeHhO1bVquIZsEFrtLy0H7qVksrUKl+h8ip27SCWbVJePwgUKRnmHysKddNd0A/+qCv477GuGaGU
AarTIT9F6IFFFbQfqXO/gXhYPoCenNVb5kZTePLsnIg5YrAC4SH+Ag6ClHtTeGNnjdxPEZPb/5EF
nmzNEDweyH7z3aJ9e2YGVNHsqyPQ/xu5Oyb1P2sOREx3/KwqIjyplXP95UZ37AksvW5aBpkgmBwi
Wttpk6W46vnWGMfL3BLO5dSa+Wt8/Lw/8SdpslVoZBxLZIbv1bqlNbAWc6S7grD2UCTzxFFh6iLF
NuFzmlXRR5oNR3nFgwTssespI4sdL84ZrOpVJmuFXfjyGVL8ue/kNVZUOoldSTN+ZcH69rOwRLxU
ahrutntE/dLiQDP1o39W6Qr4/YVd0CWnmyn6oiddq2/J0WNq5kRqriCAeABhfrj0+i1d+Sm5L7Ee
CCaZNbPAEGoEnp9v3XwOiHn03MDFjPWkncFBBe/2hWVaYslWG7/GSQ0xQ2lhpkyMwG1XaN9DfHlR
eSCbm59UzxXPBODR4heiLXv3vKeH24y7kncvReDehLo4TXCfRG7eb5n6fGaluMlZH4nJR+Dwf3/S
x2yxCzPxKoXTNxh/RHUJpHq8LKj1F52gWR7RyDn1Y5e7D/pguTTRMdffwzrjvhq2kb+BweK0Su/4
XCfUqxXXaQpVcXtzxsB/5oBqYtedwkqoUFEcd8UUnLnu0Xc0vw/icsCaZOIQxnaMO/D3ikr/EvAI
dN05QLQBDh2zSuOdKa6z6o9p54MMv8YPdLekvCugRkOwribVLEC8d8ndqn8eBStsFK+Tn43uAjt0
pQyzJGrXMyi4u8jtetLX3ikbdN7xtN/pqkSjdUholSM3v+v9z2XRBdBY9vtWA8A+JKAOFfFyw7UZ
MNQXYqQwcHYQ6sfU90qNZJQvBX3gdgkTGO0yOkWhiXbCsdIhCWTvgigi71wqCV6/ZsdUgtvXLsVi
pr0b2vpCfuTUTTo+1Lvwe2q95kmNHH3peKjmE8Xuu/g/XmxQmEuAcq6oWF1xeeym3RiycBRvHLH+
mt9PzgxluDQ6i6dDUFj36jruTIlOe8xrWt9mpalzANB5s79uZr8eMnUMUDNjALw23B8nsGMD25WI
ADzJzwaAXCIbqy5C0t6B5V9t1hoXyJSah3L16+TNn2u9wIUbQH6T8cOGDxEolqoMSRwZTpEMxNZ+
wiDAlUlZYOSiiAzIG74j8nBvLF+BWL21zRFVT/DAg7m7M5WKMq/YmYKWb/MnAkKy2TKXJWmFAaei
PT3B+mrpGRznuIEVPOf3afX5rYM8chn+bEDzjzs/CxMw0X4af39x/kXqoZ4NEicXFlaZBXlJNCvd
N/fZeWFJSxAO0Lw2aA3kFFOAxQuqlq3Nz/9RLnuwuYYw0ArXKvO9302StNo5SEkcu3z4bWw8JoYV
j37XtGRGfKqYhgWhoPSptETotUeqyroY2K1EjNZbaXd42u5NVv5mR2MyKJpspNpaH0pDKw7BOiv3
mnPDrwJPVOW19aonje96apu85jlRJdwEHoqp4x71FKJGoVEENg+5fQuP3mER51YXM/kmpISVadsd
8wR5XaXCBlRRqKYaQQ/WxZq0E2zRLOqWo9RZ9KDqOdqwUdxd1xPjzUWKg9aVdLHgISMAyUDCFkyZ
WrAFpYQPgUQdrqWmh7JcpX2zGJz1PV6O48x911Og+H1FGqoKu0wg1ON8nxS5ho+6A+mYqVV7Hxze
FgF5eNDrwKHIFJgovcamFRDc9xDcGzERA5/epThSbOSfb94Gq1wafsHwdnZV+eiAq6QZNisk9pmv
9E1dQUzMABbJpajpt9jo46EOcaOANM4tLxIR7kv7t7+xtpf8S4XV576IZFHaConll8Blw86/6G2J
v0TTNbJBPoo5V/SlCU8JM2SwpZMgLpY/Gxzhzh3bLmOXgyxbdv6XPalZKvtDxmwDD3WLpVB3g9WT
vBOMqV4sZmX9AAmcrXI4oQIKPH2trnr3re2KbY3A64hVBg4HNC/Mq8BMrDUwLCfMhZG54eaL2es5
Thi0l4kC0KrHd5LSwZrk4srHth3uDWTtHcOecewhfgcI8WZY3Qlk64X7d3i+sVSR5tFinnQZU9yp
N/f3On/eKCoOSZCqHNJP2mtBKAq8ageMetIzvu7g944mX62to+4nsBHcLzkdhKHqoAMqGZVfVv0l
XJnQoeZRsKUxFjwM56mvD9sNnXNOBrqnYoAFTiV0H//IgbxjeQcVzPAOExQ+PZUW3GCswKBOijBY
4ez8p19pz26n9t58oI95f92uZQ0aq6NmTECPZVitWrog4aGYx/ny938xP1cw2nZumgClyP8eSu2s
jXjynZSHVGdkWEeZ5uKgEO1HOD5Ge9l2QX73/0jtnnoVg9rjRUzwVdcQwq5WUzmVbl9aLzQ6KY/U
8tcSgTVSkEgKFb84StqOGicXhSKE9lerDpy/2ka4Qm1TeXiitIfYwjoUa4ROM9sWD71j1eshQ8mN
BH4I70CVV8AcLew6qVUQe5QNJ7wHwDE3zSTaBlTiKJ3baZ0EPv6l2cOvIYqzGlZ26X0GRI0GtA/W
ilnZ/aaCM/lXpRszPNJ2uqgrWxByVu7GhV3DhC23/UQKsJ7YpcPO5u4vtI1+1TgTs8/I/FyNGaza
+G4CN+4BM8ZTw4I9x6fvEIXvWGIeMQhqGA8y1ZOnF+TkVsIWhKNrpgc8btSLHpkHvoF5E9oNgie8
Eq2TYMSGmoAO9WQrHxpXgcUUUE7fz1f0oq8Bi/NWBMloxIySj2WKpXVNYCt5OaL3Qpmz8il1Mi5A
L3PF6aPnZlvFfBxlwCpPzJpWybBM7FoioRgJ4wNLh3RLe0kEdd60nKO8hsJ8BKiLw3jGXQkhB6zx
e8puxJzBs4vpTGx4A3XuA/JmtNAO/UUAq5iCIuOqjiHshMB317Ix1fJ1LFL5z75/thgq5GkNsPPW
T2CsX4cOeN8sQzsho95REb051fsd/yLnnpAF+Xpca7vvSEna03fVwqCkRNt5ykW7a4LIgURVbGkx
B7jADulb1QUrD4ItSxjCTmD6Xt2xUpjdVDRoOvy2ufhjhfR7fAdgKMeYrAIQ5luaUN5yUWdVIpWC
gyGFnXL9zqT+4/wAiUyEZUFPR8InaWPyimqfwasSvBvsj8I6mT2iMTojh3jvxeZpcPx31kTNjlKg
HcB/qffPI1dx1aViiYGuLSyn3eW9gm77bDZMuwl6TCqm3cL8DMDcY8ZCV9GGHfWrTpGTsUL+xx5d
TqtZk8rWVA6AVmuaYh8BXUFjEwu/Zn4R9RkUMCh2IntBjoGPu9x4kbu+R1XwX+UCwW5hsOHQnhu/
N6g2i5Oc+0GqVFR1+veZO2z2CbcxJVWPEzZX7ZPD7WhJRCADVoUArDcmrWu72aUXPkdDJdX3hNa5
9Yn336PKmytGEmu89Ila2AX/2Kmbby4zDdj21vafbxPtg6uk9FAseKfkOovhLpFsWfkuGkeZbhPi
lcpIgwzgpaC1yzVPh/GlHcdHCzxODIpH9IqjXkkCdRLrZZwJCCQxllmgzCvyAzvGXx2ObewK3fqs
pShvElGt1UL0qTwMGVCIJ3sBB3r8D+7AbPpeV8f0qfUNy3EVxn8L7S+NJIhebVRnRAu1bfXiwX8k
Vy6RrEYxwOmYgcqIBB7of3MhuRMz2Z1Cefkinc1X2Aw1zp2RAEjSNzkFNZaJAxfiVEaEWZ6KHNxA
GtGIPqp1ZLfQjKJgCwK6UoBCmQyrzkomjqiFv++uMV+1XGTnpK3juh0DRq4zIfny3/gHi8mxkAJx
b9djE5oLy7PNc+GB1D9tdZJdg9WK2pRlHqS/f3Wg5sxBvfj71YrF/J9qA4XS+vJt65AheSsFMWf9
9w/yg+lb3d+LbCybE7cwUAJ6ClFV63yorw6Izq7WUQ7LPefBqjbMVQELpJnvqbFGSmtJ/c1Ne3DH
9yvDKo9FaLYJkBvaIIMaDm20nB2BeX/0eSJ36q7DPMLpxNdYcrm0yDM5Stt9qQbG5mBewG+TgNoe
4jB/DKQSlmw/ZqTfg7ucMq+adTwhqxG0OTj0HWf2e8Lz6+aEFlJwLjBHWD9CYtdSfZ2ISeIcJdRL
SJzaeEHQ2u1wNz2rPTk4Qe0fprlH9tu7KlR//FRhglpcZBR2qAfZatrOdFwJFV+saxJXNv19Ml5O
Rhv+MhrsfbTKdbbh9TnRRpWLhTuXIvIlZUHyyv6s991hFhErPGqddweRu1LfKru/k6WgEh9Cg5Ff
6w7Kw9RDZ8tjaQDbfIrD+U1eTsONUEVevbaRLhcYX/iJ85KwpMic0TWB82s9fjWmzwimEnMO2E4X
gkhyU4b7LK3eLdrhJ0+qbQl0l9uygmErWaYDNI9WWor0pQEnC6W/6//Eo3OxcgQtxyakORV7QqxH
5EpB/v4iNCTClj556x2iW+riNfAHqgmXjFLOUKUvC5OUzvlPpchTfd5G6KLHpHDG0y085QYTLHe7
5bSKHw+i2s2eoaiGtzEdPKWZ7S1AbLJY+zap6yvAyFZMRAeqZJdx4eM1N0iCWtVM1lchtUQa2Hgm
LyMXv9xufP/OOHe8K40vvSL5rQ/KFVrPG9KqYl5jfP/wXXkG7pOxzdk4Fle1BiZZLV0DWgd2sP7O
GKIFw28HwwU9q1ghVjXQoalHEq9nvFqFyc07elYyomyMm+XD2WUGN+fkIBe/fj6EKMwjEE934WMM
tKCaOzkiFiKAoq5yvm+3O1TtpQH/O1DwyNM9EAM0b0dLKCz0dBqUrPkSu/M4+CHNtuH/DXvG+YBd
Y9TWeOBh3h9m3pBB/KhQp224Ymdj6RoErtKbB5RVw1/XpmtaYq40gnXPK4ERpHDO5XY0qHucID1t
Xyc2Bn6+HDnIV7qHf0Ma1FGd1KzHJ/lBXy1sny45pcd5H+iA9216KetsJYkVXwORgw8AlnlAWBzS
6NE9wPsYR+ekvPiPO7R3AkhTPEKCDTTR1NfMQAFzBKFfdnmgM+j630wMcziqNwe/9YT4qEKlv0Ng
1ZWAv8hb51yl+M78LRbXroYy/Mc1tO+p9uWhLZGA/GTLsra/ScfK6W9k0VetdP69O0qLGz2ehvlN
5/uShyeyrV9sRpLXXrBFbkahCNo7/Sckndfm+l8r/aIxyRoZuurgeZ8bG5itOrRf6xZzo9jw42fN
2r3USxSo1+XPsDCjz7bLvWQ3BoJkZCw49nmC9TRRpV+S7pD4g9e46jqFpXqMRUI1bwMJWpjW8UOa
GH7z6SxePg6fPLgzcrH1rcV22brXqBSKXtfqgvX55TC+fCev8kbCe9FoCa8RAcew5TJByPUC889r
4gZAxYH7XlfO9BISsWz75ImEYaASZZ1wRoADJGl2dCi+T+29PMZ+3F/+sdtCrLWOjDTC2qibjrYQ
wBbr0FSaqM81WUp7YNszCco+JPV6tlOouCokRUFTaNvD8tVVebjC5oRB4iniVAFy+VgUazXgH3B/
gpB5vhnwnfLCEAWEmcuIxV+/FN7Cj7odvtLv2cqzQpi5xwVVaFl1fVyaZonY1fygomIaQRLv0NQv
HWeHjfazR9lDJJyO61dGxGcJl65n40vSLd8Dd/vdxzPQB6rXE8lxVeB6x4S/MhfsekGH0eCWrvbB
UzH15aeUfXScmZJ+RxrTFkbmaLrwIdJaygjSalrZjH/WXcyt4oIbczaoOh+oL8gGswFRQUCV+Cgu
XrUg3hv/18PfjIchqq0vsgpGlAQu6MgbD9haliSj6R771Ke+PN98HsRZfwZMnPXnyjT6AAUyXiwo
laJPChHKgFpfddGPzetP/drfy9C8DxZWRwOXS4sNVYclD8/luWK0TQu3jQWLzqORE+LdykL/ZumU
lBf9eaw4G5nasYa4Nv7DOOL7MdPeL4H3U5n7xMgordT8pKxpbLUOeYtysHGoMc1yn45PfBZnhKUq
yS3eTYqPYseSrh+qXahrh344WOk/V+RIM188uQyQcH/7HtsCCKb4SJHlItDvTkKGMqcka2ZWZgAG
VNyc3fU0/AYz+fj+u2oNZTKteqSruonFcVioylhEnsgGChJ90ehV8fU5iE20pvc7vgZdkrCWsg60
2LsJNDP9bOGF5Y3c/HCa6uMeo94hjB55MmRaupOhXeQvI/BurpNXD9P3eqCOuXuPfhZn3OSWS3Ak
JmUe6Fe+ZdbFFX5rUxOoWAF753GxyJQMy/BmuMPzDeD4wgYBP4Izo8pFOifjmZz3Fch4EqhEECGC
Aco4SpmPvc+W5gTReFEGmGFgSUE+gC3dO9m8h0Nq4D+gVuew7ya7onjIJE2lItkcbYmiS1GKXgXZ
dEvTlsYSopfToIMoeBNmpPSvCB5Xs8coEVOmlTV3XSx5evc+lAaKcfu0hRqN+MSJ4QqpB/VXwS+a
bL6JfRc+CA8PCWLQgL8cbpeubEKJL1wYtKMsYULRLLtPIy9oOEBy7sd9+YsQDaetjnKAXIRCvisF
x+33r1AYT3OKomlbpZhNrKnDWeYyDegIrszvx24FeApsS7crJKRumecg53Im9uUG1xeHlDqAoiQN
qBIzmPTjPIg+JMOGdnf7Jed3glTMv5cgr5O/NnxAFWj9YHymErhWJoxtXcN43nGaA7wJz+poAjD5
UYhmdFkxZfv0KJmnLGd2/Iu+zfMeU08syzp+vosGOgAMisZD10o0vh46cVyAmipICGCTal+60wX+
FQ3kyFPXxGM6Xs09G1UUHjUfDkWvfxLbgMbZKgpcHTQPTsEx4SO4VJ8DzwDqjXSvjMVSTX7QuD7l
ayu4bQQZyKNPy+/rsFDtIUz4C+JqkHalSjDDm/gInZL1bDLUSEBdAS1JZelUTNb0arC8et0drT4x
JqZLKNcEXE8FeDcqJTUEFRQ8ootkAD+WuMqLZsGVJYBaA2Gtv27Hf68jjPVUoCqmHY1MAO5nna8E
KPyBu66neC72w9VK/YvXN/GtP8yjyiHjr+xhl0HN5z/S37QHNmJLQrPPnRkAE51zZTEDgcaTp9GF
9xDRE+x4xEqwjzXPYxO3Xiv18jKW6r/bFFUYFcJhgGWCYH1Ug8LaL092qcTxdYDDefihUQN8jydD
pUFMtfXivWEwNEcbH37v0dSnxPGite5SyN7WYUoIAYa9cGHdU1EJzEjwNIovsSQUsm16+hGkKTLK
ObTzt7Iv9OCaQMQu/sjW3c5eRsm8sRcbYOoKDAKbNuM3ahod/Zx2WmpGxeTeAZcOePow+TtNbqXW
Bmb6PA0FbA575vr4VJZV69qgU2dj54e1XEYut7K4IA8I/Hjvt1g1s2ytWyo9pVNtBTZZuTRl4Hds
ZRhKp1AoXZ4ZkqR6oiiWCSrkAnBPDZ/8AT1BoEbNYCgVsfOp3wBM47NEZKRvaRqGzZ3LULkLw8FD
vuXOrmh3wq6zPcgGKZatR4wBcRb2osJCEgKTqugyTRwptxai0SvRMn+tuRbg18ZQH191scrQBt7K
CGSmCNuPm9Srw0ia3qnD6AAKh01jBr8ct0kx10eJkigm13n+OkDeqfW9xJpzWNocXlDbYoeU8V16
7NWT9Z4/aMlEzgCfdLzomhj2mV1bDLTnfd7D3RFpcr+7HVRm2LWxNT0rD9zCP9BdJRrILuX4HxuY
8oBfbEb61K34vJVOnfXxI4YIRYD2CxRMFohB4e0/GBit/TdmzhFI0L3b6UivT1X89UsMnR2oFBig
+4c0XFCUjwbGxx+LMrUOWK0COwLHjqUtk51p87Tu2FBChfPfdoB1mJK09yXhbZwEo8pBUkX1xCW0
5/75UwS97/79QF9MFmhiCmTQtWalUsfqjQRvUwQ9GpHZCTFD651HyPnRxUwjR8syKWLj3+S83kUS
dnBRknIZ18gt3rzLrEFjkcileXcOlXCLzyph5pVKvQV/FTgRkI6nc77TuLwvRwegehyZ4pk9Sevw
/cIhpaU+uTwT4vyFd3M5z6HJ+su66qa4S7E7U+I/I4L4wKkwYa5BBW5hSk1WVaESb5ywAvXHAd+c
+AJWHw/lxsZiuoMcOOVbUMxiBmNj7xhvnDItEPjZcoKbKiCqZvTp60JmaZGxky7SYwcYG3hEAhaj
iC1zUNSZvFfA/SKVGhHgfHNhPp+OZ0a+DBfE6OakCbGkrWJLlfyAudg3ExSFP8PKvFqVDD3qeSE6
gq2F+tisK8yqlkWnIlvqMhd63+B6jalM75TXX43hk0xLQH7aiz/Wmth/r8DvT/l7RUfDqJG6LYHT
1ZkHuUq57wkk/EikKffyyQgkKXpgQ+DpvKtcmKeJQWqKT7YYXvf7jVN8afULS9ZQwhOigG0rcKjQ
VAFI5OdPCYNiqDGANLyXqqfX4sicKBKRb+qrD8KC3VJ4RSxCihFmHnlHpc7/7dUO75Xcx9yCNkxC
9jCWzqYkNf6Yddln88QB28UM1ySi0bpiNRir3vFnD2Osc/95vcJ2TRIFm626SJt0rF8AZUcCX1Y+
skVqvcKSKcg2rTckaTYigoQ7AM3VuNdyQbG2/TPpRqdG+B/InyBCoQ+/OOnwXUvBx4SXxB1+8VzQ
oBxINW4OIMnEpTBcD37JaikrtxX3fxUjY4sj4/snXcw7rSELGsKpaEOgYIslpK6SAN580rNl/+ad
bBhU30u7jjvdeSOuVdyEq+iD0pM1SWZqEc7ceGbdBpCuHoBXqk+s+F7qiKjK7ykbP+sfn4Uqlqi0
BPbWOZCwpHShH8GkZhpAPJopYdVH52slcnFbnakUR9E8PZIy7j8SSAzwYeg1FE3hDwbrbBDdAvL7
IBq+/1br18hZ8f/quVCEIhzG9OQuXmMfTSPiRBz8VjXn37vvV5e94IFai/plQ0dRXuc6e5cR8yTS
HJQ6La17suF//+vCeVDWzqbwRh4kLeB5ZMVIFzoFOYEM+Aw5ybgEBYFZQ5iooGzhLtWAg1OPm0y/
htsVqNZSopE/ENlAh1DHtnkMDalGRei8YhvaCKWhBAruThwgR6bx8Eyy9TyvSZe97CefPV16YA1+
hjnjNi4VFqcfvk9vYzUujM4VbZFX9P93neJ2RrykaBjC+5u/m7+HWz+vce2xy8XcNFJfzrhHy8w/
EVaetYSEFaxG9rkixd1JoeGa6kYSSK0WR8jhbfKk9s1wsjMcVafAvEoxNCgH/L+qvbrtrTuu3gbw
eTgBaHp+cVlAH9Pz7HYZD26FjKIvePmT0+0X4owC0BymdySZGRwEx9X7u5j384lZx7yfmky/Qazo
6LK+d+cVS1Jo3z1tTG2q8dRJnw1yBOb0/2fxq3xeTjkNXKyEj9z8/h2lrbKMg0Q9bPrlUIGb0kqV
NZaJ9lCac7DqoO6+N8zzHz6mthUpw1hZpaCsDPBRcB7+FUQZjMxXVWD60518GyqXOHO5F7XgeIhC
yMB96ymVsUsEEx56lAfkYR8WKvdt/Z5Qs2e2l9u9IYkVGy/uz+ov1eYNeo5MZ9Ef+UkHtZ98Lyuu
/A/GJtXZ0KZDEKU7cAvbxlr8jvG7HXGbPY/GutbFYLjShh07ycoIU9yvk9pIQIwwHse7NDyBDjow
rwDiEdGkiITDYpjPiEqCL54zNaOvXdVrr5mPH1T2gvcnK9zrP2hcKBMto0Fzr6XkqSBoxmKtxBdU
qchnhX6PRx0EftZLdl92sGqHpsJMyF3w6EThICrYbllAlRbopbq3aVHBphBpN6ConY02M9KVKSA0
r/rDlAfWEOpELfikELYO2zLb+hRpE00+Tn8FZxrtaLZCm8zFr8P8ntRKrXr28Gs92fyTnEeHveFP
D0uykFJwBIOdc/KnWOdxaY+hv5e2VSMU8i2RZccm85zzCqeIpw8C/0xoXGeR1LYV9j99IKG4br3C
UdQR3Eb4ALYYIWLix27shwYTtAOCUnQYmy0nhaxY1Z2cVjeoQ7aaR1UcBTWiSDMmMW8tArDGyEJ5
fd70fRaqPbBmJjewu5jhijMwG2f95OyWdPL2R7x4/E1gOCd+pu5954vFPiIx7/FP627SOiRtPsZ7
L49P2imZEOhIJGLwX0n9iuIWcW++LFxdiss6G7nF/MYluo7nytaXUJduyWtLB3EL1AbxastcJ8A4
krQgCUbB0OAQJLfAJpBQQ9yC3BYm+TIjITIhGAPRdG4JHYfUKMqGyMoOZvnqLz5fDIbk4sZlTGU+
M9FL3b+02ToxFQymkswKdIBjoHC7y6Wgbww68G3k0OSYn8Ry5OuFntHvOWb2p2pXTdlwijIYcok/
RPPeCLb9ljA9kfev5J8+pIV6WoWeUBClPOwosr1OwyQivur3GtJXeu/cxuSsQbeVuVDvYJ2GU/Ua
iPbFqUMrxqSUzIX/XV7ARILpWPHK5sk+HzlHPESo9bOTiHFWiG9garmkPZULuYciyBrXXj41L1sR
myMqdvBkrBS5mA0pRWbJaODdp4xXtS5TrNIDaNtMM+EbepyylfXx6q8FENP1sNlwRIYJK8j6nZzU
oNcIq4DZFaeRIntKBxEQQ5vMoOxcStDo7kpq2NYdSNcrHHmY8kraazlMbRuzakuOTbCwmaLr7aM9
bmVDKM+opv2W/akEzkm3Z7MqnF9+z4hvxPcl3j88jGNBbLmYIatXCP15iC5FA+h3G+nS3Iph4yQu
Bl6jlsIjC5GBLC89peEhkqZ0xyQYPsK125AxyPQpw8xFhdYi+gAk5ZHIxwtDe+lHJBIzOBv7YsCn
pHL8+0boRMjzjrvoP4bW/fZUFfvbxYixZERj3Zrx7ElPTexuMB+0uSa5rYw6vgOFfcREIuAyEXzB
V750YrO5TXNlwrwmkrfp76ZGRHr989Mc9Lk6Y/QoGyVnnHDb3cYnbh2vEV7eE63quJlz9E+yuyTO
8LpX2yMtkM4KiKq48w+JaacwNUaHBxHa3qPzMsJqRRT19bKjmzNHmr22Y6tZCWwIorsVPbO3BoRH
oY3uySaoJJJXmBoL3XK0fHI8QW8Y0GIGsklkHDG2Mk8uDTnpi6HQXT1E+G+PQt+WQz/IJssOjSYj
shT4B6lVHIrAfn6Ggt689aN3YPP8Zb/xDM9K9xmc/QOwxHDY3ALyK0965hE2L9PDpgH5pqVNETaG
jP6VnCzzmPS6JevV4RbFKfYMAstF9L8hS5KvcI47r1MhQeUOx6R7whSLJZ8mUIjUkAsQGxldbtEK
uEYc1kKbim5/DvtC3ufVeFn2k38uLoOkwzoBoZALLHL2RqgWRp+Gd4tLGzvzmX6F/HqgcBj60ZEh
rp8WwlheR2/qN5RCY0d7yt8yLB/XNzCrtk9xHlM6QLxRpTYol3LxwC5w7hWqur3XWzAJ7/MkqzPB
LKx11Gjq7wy2z+2FGkBSu/jtMp3hqsCEFMnUdpUmJnKrrTxvIabP2amQBRvmlF17mxWgRDBMFzMv
zekO5ARAe0FXiEwy9ecUzgA02SsGI6Rv2TLgkYEDTfgsLsxS9BfVJK+e7mO6Ao4Z2BijAxWI/iGD
9sr+fNlGYiMPQPLHYJ4byp/kw/yULNAcri4BvkpaxRlcnEV+YYMRIdGlhh3oPjxQC1GAj24qGE1N
SCgI2W3LOIC2TBXqr6rRWW3jogoe7X83I2EgmL3BfXx9M4bwR+iEebIo9TvbellJOMikXCyuEk6j
n2tcmLMUSScWJppSZn61mPLsMfqleMmln7UHLUYIEHkmzDu4e7m7ggF2fK1I1FCoQ4f23QT6+XVy
fvSLrLKjCOIEUNDdmxU8frjQRIZalfvJncywefJoTPbQ8Lx+nW17NsCjPp+EF0SNjxNnHik3X+UE
bd9y4vkXPbT34n6RPgzPc8R2a8CkY9AzaFhfmyF1+GIU2lLDmEmEbCPuhrxiZo9cA5AA/7wKdbAT
2zEn8nxQH6Fjkmt9V/us3eoKIGPw75tDuV0+3jBxxYlY2ybRYgOGgyJCZSDAHmbGWxV7Bpv3Sz/Y
/Ob+OytWV3BinpyerOWFoZnv5N+yo0n3S+K0pvQcjqAZwIUlft5Mw+9TtrGAeRWuFB2MejyfGiLo
sDVSkASPbC3RKFJLUA0NA9X5qi1GxjJsiTB7KR7mu7GSJx6WGacgf1+W3tehZpfoFo1368gjEyo8
sqHA8KDbhOeibLnAxGnXBOnOue5591861zAZbZWHZKesRRWEPaxL+h7uNgu92eIIjmSpZdwX13Bn
k1mIcJG7/PGN39Ju8H2dzgUN3lwpnZXgJodXZOc9as79Zr+EQc5OG7KQO/WW+potj9NZIKtoZZh5
VroTUbYmy63ScGmyh3cmTsKbU1x/095koj5HV0oPoM+EIUHzYAgsG44WH8xpqHtN2q9pFaVn3lqr
42f+rLETsLYL/ZxFvTsYfUD3QSp/TC2v/pV4Sr1VXp5bgVO9ZcA90/PA4llO7gPvRUFuyWb6boRS
sLp58LnnEerehkBmiAL96j7MDBlMzpU7d05S1UWC5oU82zPjSjXBRSqx10lBVNuCQN0p4C/sxSzj
4X3bOYH4oTOZS1QP1E7An/S2iKLDxTaC5zQ78QuNGM3lPbpPLS4cfzLJrJUp5F7tj2ZNkZ/XtYQi
yv2/pntwa0A2N0r1GWdlnbHTpJTtY9DMedqp1nhfPf7E4BXwLEwSomnqIB19/Hh7Gf1I5kR6or3T
Y13Jx+jKf/SgVj0xataFi1d0n1xOV4eW3VbcEQs+tR7nomlvEVl1vbMsPF5D6dBLrrKnz8N4+sHA
C6wnJehpf22t/2hGIzE+5hviVAsTQmtwdkHjUR08Awln+bxkzFtcRTD+EZoJp85UpsUXsAdlZizB
hMiP2/BdKf5YxMFqwGpPCKUsQ+p8YylpZOKpwuCfZh19UhQWlMUPtGyIjHNmpdXmtxWWp7bSPhJk
06BQqIL85a1h8a65/5wrgwloy9Ztj8z6qqBLLeg+kG3ep3N2l9n+OCSRU/cM+Gi/xNk6GVMZxU33
hxpbQpuZPh1XFU/Lk4pjcD9LQD6w9CCpwjWZwWF/K+wCxRHEdvr5rO0HsVJZZj/J9BE2G7OVeX8s
GYfsR+0wRB4TIyRY7RGYLoi0srytt3nkQ3dKAlvZMCtIon05y9f7tf3gDDQBzFuYqUDufgvooGNE
yxBEqkHXaCvkzG/ECh5No6GMRrgJpv8D5hQY3bV4v3669HwsbwsGzBPKqRpJIFG1glefo5AEQ7Bc
d5+Wttalla8BSjW2eLEcgtQkK9gbOwUi1XE5+rfHe1N3QIJk6z05L6mAqKc9+KfzP9qbD6YnztGp
KhIbSZqimlYCDcVvthz9Q6ghN/vAqNd+FL5xmkUoulmNa+l7lobLJbL/WquWG8cCyro9O7BD5gSZ
aeZHQ+LqOGJ0nCSQsbZu1nm3MHh8PSgEOOiz6VR2mOWgleOMZLuFc95PVA7yteDmZ5SzOycFaw8a
2Se54xz1iOJO6xPpC+awiPyxhsbycxd0o/jR9inwT+Aaq+IgP/7H82k/FD0ZW/ION4EgmAYuPp5m
/GvyJkhKmi+CnCMwmB4GLujeck6Gb18sPAMIt/FKGcxZciqWj4bu4o6F2kCdWzT2QRvHm6tFzclp
6SWsYBks651g4f8U2Q47j7z+oHLYq+XdSq+9N85f3ZHy5/IynOIy+Rwx6fkoU/F73nX8d1TRkFeV
1CUeuD/MvuhHoRNf/Sro2enXozR2L93HrTX4eG+wFOmuv5LbCG0VXy4cHvz66UKTwhejDFZ8GzsE
CbN7lw5E7RNmLUb0MByvGMaqsk1CGsgHV2ZQ/6yqK+ftau08AmQbd4fZL9tHmm4VzCM17fj1VRNQ
hEdjb6/VGNYkrguj1ZtZnOXdYcLQPo6dR2TCx+VVJ2GsyPoogk32/+hpmAC3Z27+14TIp6WEvNOR
HW6V9N2ljyFa7r9BrCK8G+jqRFvA79pb6FW+oEyT+Y5/+xzxksLXbYn+MysyBM+MUwr1gRaNem1y
gB1vKOL+M3fh8yFIVmHTXSNzxIB4Qzk2BT7VlMUSpJ8J16I3vT50lvrLagWOfwZ04phs2wl1WB3L
xs9FKQ+E60q+2F/98XbQGOSpUK5KH1/LPEhDrCeONBqqN0k3kf3Qj6j+Uu8/h1Tcfbe6HI4IIVoo
R6vLO2IC7sUadgtRv/Nfnh86twXBTxlQrl+TCulsXDooGAUNWPPHRh//bKCKfzDaFuYU/F54kT07
Mm/68AamOF7zqQDW+mUOS8vLPU0/iz2V6FIc4U85qs/PWr9cGWx6AgqnSOSBVXAA2Qcz12p9swjy
a25beeEAH87bu+MOFsEQl4FjFLXhSdNWXw2TrcOWCV+HvSXB497JiVP+9PLRAHBXkRuKk3EtC1mt
XAKZ1NTkqF/hiYQ4EFe2soBSBho4FKmVj8WWTunxuIDnHzuuOxTLluw+uInyGZ2AUCItbmce1phw
srolZiBYx2+PrM9Lm9zcaFXwAuZBCK5hzabTqV7W/KGBBqdad8BB0XwlCti7xVtXSJSHEATodo8H
92/ol8X85/Wr4hhr056vDTV4XB8B3nUc3YDI0fHv3C55Sf2YleDW+vyZWgTAPYcp05RmM6yTDk+P
BgyG1qE6tQRI70WGw4TH9wNtzRvR7L1hDCW6qOE2RC9ai6foDU3T07TrYWYbBeu4D1KOn7C9BGXU
U8/06xspmFi05XFTg0JS7f/h5zwK+pienCFWUoCJwDSWj4c9apsUqNMylDixZfm9/2fmixbDvFME
QLOBTL9V95vABEiY2ub2Y1ihaPt7Hn9CBEfBPE6PCmIemWRtLGDADbewFMVY8bWolDkiui2Kjyaa
TPg/kMlzPHG6hST/Q2z0+0Non8c1Epoo39+vWEp5BsfVXAel1i0DZH7/xr4XikVb5r1wv+NqUj9U
cLJ2dIvc95P0YGWB1/cQqKjx0WWFAVYcja8bbOmDqsCrdPanhrgOBo7EEXNDREx2PDEAt0v8A0fH
l1FmPyYlf56nhC3wPoMtF/vE9sKKXKk9Wvwx1oHUiILs5N05KTlJMOddZzrqWyate0kKkxGRogq+
AQxI94rfLjU1j49ay4AzmPiBYivn3GPa6lNsE7CCa08j7Z56iWKMrBNI4JQOg+sWBqa9q/YB9uRQ
yyNan8TgooTtap9YjAITGlpbfvXtIObCfzTSPISf6sZyvGR/adw5QHj90bxmtKMa4HBAGEOhQ4/t
Q+C4EAorqnZtKTjDK9m3OOaJ17ixHns4RFdHKJIWXfZQfj0Xu2RTc8yyu67FQQg0ubLXD52FGG5A
k4tRqnpMYO6zKEVzqgBKRGmsnANhuONESTM5aFJa7uTU6FiQ9q8qipHMx4Am8tvudcJ+N740IR/t
gaWrAd/Ii3L0tMFMxV+HDt8Y7t+Cw1bOXpsTWe3N/QlINAtuy6RuJi3p5wt8Z+yIaQLcn/gYE8LX
J+u0RmSaXUBxZH53C84LzWTDTKpVvxrAavyZvAboD96yJah93bT/YxdUAHTmnDS2kB95hM7Uuhqg
UqJUypR7nqEdjZ/MOfGuSJpJXIQzr3LUE5QaFs2U1E9Qm2GJCyfCv1IUYbq337lC/HzziH815fro
saXVv3crrIRwhB8sS/u2BVMCYOuvpsSdgflyVbbaeeii3tEGxOn/xjLJXRue0XTSSdL6enAojuww
If5CUjct5lLGdlf3qZNfYZMI8zke5qFChbKT225Y8e2GK2PTSMyy+lt2gxRlL6yhHm0Pz5Ym+giy
FCln4af3XDMhyIZ9KZgweXbweeYVHOl9yJGFoPHp7DaLzoZf1a8ixc2KwvynBlf5V7EZj2B8rHCM
3mftqK1gOHtcUNaIWlaPL6lzCvuluM+KNn/KIfUBgj0VGHzp4/P89iP4qK8gJT3Gqpzh7ugtqpJP
m5Q7oLjPYRZgeOx+kzWTzsi6lOtjP7U3LpkN5/NHBKi/3VqosFgs5n2/osVA9Q2sFdeF0D+KN180
AdqVCSuFMS5+lQ9Uhln4s7B04acWFzJ8TYZy907u/kOTXNw24o47kxRC2rmnH+ezbVcfd5idXn/n
Tuo8UWBV/sPR2DnM+gQfbT3rtbdnfy9iWrYNzoUdOcFY0QuomOZ6qytAUX7FjrQs1/4JNsB+bfhP
fUsqR3sdQph7ieGJbMzdJLZtWclZK80dePz+o4Gq6aguipufjy+FcKKkWhDjHpsZe9Pa6o5ADpt1
OLvrqtra2OaYh/RRBEcw10McjhhutE14HOrQDl7soYKOuyXJgHPoOOyA7eFErPARDrYbQW+LZihb
NBV8jrEji+wM+tgbfP32Oaxpl7IU7gwAWt5WULx4uWex2VvjFqH1PHg0/vxJ5xFbbxmHsZ2dFqGz
5bR6OnmGhVz4CrbRZLrl989e/VjqEjRkzUNRH6uZBTF/qNtNL3i0vUBiP8EON1B+QuM5TN41Kp1e
EeaHU+1XmD8eZWO3lqquF/0DLYgA1QRrIhEjaxHjuft59DQQqAv9A1wLBlsu+f4teBVYi9E5NGzk
HEw7QML+MDSjxzrvjc01eJaU3ZP/9w8JnilHsZ7WTLmzMs4a2opdYwm5J/uz6JU7PLeGG5BUue6Z
kezN7Jwa7g3OGHZdpjF6hPCkTcldmrS2JEQiAXnjCpnwFhkgILDW4uTcPeR6w7WKXkgv18+5SL+k
ZqCFPN6cCfAH30BPr+9PJwd/HXd+Z+spsQgjtT3z/zZ1cBVlgRdj0Pr1GefuVXEe3I7H8Mgs0izI
/9/NVc6I4CvEtweWhsmYIxYPXW0Z/0M7zF7uiK5FlAXvrvkYHhX9VnCTBd57ExLpNK1dlccJJQpy
1R8qrMp7zz2cZrS8uLzrUzK7xr39VJMgn9Fhhn4+BI3RVciHaxPAXU97w7+7p4OFQhyuHXwBjyQu
wYFNPPD87ERSaQsLPkPADUElKn4zmJ4lPn6XvQXxgSFuC8LtXRFKUWmte9pgP7kMmSF30n4UE8pF
jCT07JUBbS00NHY86tN2S4PNjJEYkBCxiuT0FlDklV9Vt97LKglrWcoiCUpwYAyhbWBZWLKKgSDp
/8ztZTh+oIvFhr6gxVTmOqX8LYOTdxZ2U4o0xE4EsCm3S+NrBngMM3NpjgqsV55JJRlU7dZ/uaHR
kAoxLZUi1Ggsy0Mh9vjntM3tlFu7LkvlLCit5j91Qe+Man4ammwABMkwIeQ+VG2t1ds3Ho9aFIeq
7YtsSkWEWrBphs+sw27yYjOpZO1B7q2PA4mUSKXdv1pzz+7Ln1I5fZc0qpu6JjWQ2YYyFSfImw7/
p/Jbu2yhsSEXmugnHcS7OR00xWC3bvUnt//Kk2XWMq0KuZw1Dev4i9eW0Bn7OVg/I5hjHR7FTpAI
yEHUnLsysr2C3TCUc//L9jlUxWHGTd+6U7JYfVYCjGasocXHCKsEFYUOkudBMWqcXgFmVokQFPwH
pTLftSmsyOC6Kn6aLdGsVE4Q5Lr/QnSTleLu9mHPdKabp+Gv9LjRTiurLVchONAqOsFQu52fittb
3DAUZTOqIFLMRgkBilV6kTrBr3fgCbnVRrqKGjjcbRnufTwCZKlHINEUXcbt2JuOzRzWZSaE5bNV
7mkgqKAq/ch3hI1803RwRk+W7Sq8ttlSv6dsfLmVRckdhMCaiBLfl5hmyOMBW2PIMO0nWpofD2tZ
5oR+WH8RefFkFK7JjuxZAdGJO5EcX5nsnLRReozlOuYOfyBEEizMWjyzR54d9cnNVxUTN190cEBb
7jQBAbrYX8UOFpEpVIhJMcqkSpdKihzHSM+QlwnqNlJ7IuPZBOeJioOpGtKcA1Tf7tM1YHUGEHsc
f7GeqcpGIKInEKnbj3Ycn5bMyHRrv7PTp3PfXFZtjKrt2HizztCxWjOzIP+salJf/pwtb/O9LDqQ
3kQcMNxSSPSDPieZXqsRBb6uts0CnLdXv+cq14+KNwE3Q+zkSPfbSJuATEnUwlL1gbPftrcLhuV9
3N+iKViGbm0IgKQ3Rbq85KTU3brTtu9Z3rTFaCkNQV4jcnBG0ouM2+dzVsZZvMy2qMMEi599Z4Z2
M29ZcDu+XUstvKD3NGDLnlC9BhKeF5qRqKpwVeU8CZGxxt+Hp+CH24EIEHnXpQ6m4I5sXcgwibs6
NF8Fbcf+VjaZuiSlYmk/8sbcpJDFPEumCkDMRFHh50vqcGyKG5TnC9qJzOLLPOxU+h0gaMRmFuT1
pyGFuGoxCNU1Lgm4FII47J7ubxPRggYSHgkl/QUzh2FAtbAKeox57q14+wjlZUYRSAJO5ONB1OGQ
yKYAIIj54HLQdHpx8yu9+VMmdi91pJDBq8Z3LqxqFFhKyb6Qp3F/hQpWHBPvRgw5az/4oKZUoOlB
3t9aQzw10YLV9nys26BsEAJ4zCpwXIPt6EgC4twNlDWrFM2DG1EGAbo2DG+JJONbNpr0d/8LGy7x
A0MdyMLwGH4uh7kakAV6uKujnRM++IRTEM7JzxBEG0WTaYQ3VDmdH3ItcgVxLlB4Lbi3VzRkDvkh
l3Yf6kqwWyIMGLdZSWOgFKPhQ4SPOBlFhjZhDm9W
`pragma protect end_protected

