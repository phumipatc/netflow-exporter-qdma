`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
B0iaJAq4pozO5ygZKBU7ivhPr6SmllDy36iovTc8xBtBPEb/197lth9TCGiyO9+5zOlBCbHgFDIW
b9c2CdqfPJ7JoPi+t0MEi6pD4I/nUQEaKxg/t3fcizY8wg0ShhxNh7wEXPI0osFaga/Ga7RPd8jP
Vl/9RYffx25oRm6dPwh1KvzNB+5WHZtzDhAplPISuQgImRzhBvlv3BE6FWLjV7go0Kuwu/P8QVnN
WD3N9YKjg9K/1ZSEyt86VmNr1OoyFyUO6QaH8hXk2/DOm6lzSEeI2GVda2XLXufTj9x8lT2yyUP8
ryEfY9sNL7/dHwzBvK7mec8FB5+K/nXtLhNm+g==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
S7+nzy++DakXrgoHCmSQpON1g0SrsEejqn3n+uk1BJSBzos2x00Yd3x1c19PCDyqvpQLQvxNYtFs
OcrE5odxjis9y70+biPq0/Yr534Mi3Ymmzgwq/xmRGI5vOqMkBHj5MUnT7yD4oyZWtzxu+9NPqsY
Ivqma9NGrV3HlMfIwXnU4DHC8EVlBZSV/JtL8NqIB62ZIXk/yiKB0g84vRgq1QYCDOugjKY+Q187
e1AXonPpztfdbk4RTV7KB5ciA1jUJ+IjH6sI8dFWyDHxSjh1ka7jDOdRVVkjCTRokgEDWfcCLvQV
SARk1vDywyis37tQubYox5MrRz6Y9YYAvyy4uAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
XA0rnoiTzxj6W++zKHMr/BnicY3bIl99eur1WUXcgNCsIBSRKAITr4u5QTclDGn+DYlcY7Xn64bT
5L0jB2OXvw==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
N3Z9mEEImUt9riHl7PSVacZJJMuNrN3113IHrRuddsFcuCSOVszECd6w9Lsiw8htncWpPBBbbfjC
yJDUKY7p9bhWA/SqycSCfRP4mPdFfH6sNEkmw+2ijaqMt+y2XspJgl8xcpUalfqocX9fV0+0HbsK
fVfD4IZPXxI23bDEtfjNK4PSCPACwg8mYH2Edvcuagf4D454ZqsocRGy2PAH1I1FCva3yguXSzRg
9yR/o6DOWot41DOi/EAkS9SEg8VgF8yvjUrOWJL83PhtYRxCmqL1qqVxdhiKjGsJI/wk4+lhvZ/V
h8L/XHsvUYiLcQS8vNwtGqtNMsL9zWz53FRSEw==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
iop4WuJMeI+7y2RjqvY0LMug7SCzEr6RIXYffoZL7ZDEUov1OU/OwrB/6Apky9noGxtcS8K0dxsX
vCFrge5XcRFK1prgTC6fnHN8ZN766JsO7JwCrT/Q4UZDJXUMV+H32+q1KeyniKFTu6JBnlWZtWxK
Vy1+ygOFqgNX3KW+pKlinoLoG/6qAAQryAtG+dlYxRI5bAdRuxkYA/Lsn+Vmr4FcMs79MO48LsDz
q0/0AJo2ntczvxRIVin+pEfCg17YmOYm+PxKmxkz+dghs22SaB0vU3ix0qcI9Uj1HxZPiTgdGvnJ
aVGzJ0+P7Rdxx+6bO61115+q0MU3ijMlwFCS7w==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
D1UpeSipFR1qXR0xevmG+Rlqkpr90tOCLEfRtk3vaYClDNkX+7RF/BbY+pftVpfiH6NorE/8JwIm
qV6i0GXe1Qm3jrpP5sWUOSkTqAZHiHwuey583gbVUys6DTi8xv4eYuhU+D8ZewsXnBOQwadlJ5/u
Ex1TzkYyznPYeBy0G3Y=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ruvgz23+J1padP7YVvvG0fwZk1HxJUdyTnPt2cyTHrIGMXxR+39g2uyPiHPkocb+kTLr/QtZDFyh
RValGCXgxZVJRTRrAJJYTWNZIPOaMk8A6UYk+4GcP//8KWU+Ostqs0CfCw1pLTWqEIE+Njg7HoqW
29gVEecS9d7LgJhKa8Y7lfXz9K84BTSUibDS2/ux8I7SSvfeapsfFHolvi0CUmIuESOs7TbGR5ga
PfeYBYd7VqEKRPYpq1C2m8KWPGwDOvXHWRP55SEnBSriUu8XHuDOclXL89AYm0xwV35xjRLV+6Dc
EUQWRIDOCuo8l3X+f4dzcH/0AjD+y30j4PxseQ==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ys6XJnJ7ZAc+zOtyqpB3dGG+gLneitnpU4XqB5Om1MLpnMDNOQ9ceBL03esWSpznr+j8ArrffQ6I
DO58Bx//apJ6ceE3NBNK8Y2B7DXFihLPrxj8APUvqoglDE8U0viHqO0WQMIHaTXWAsjyUDL74Cqq
E4dP2X6d4IzrXj1Kj7lrr+bL2vSW3QXwHtAda++XCI5QYu/Mtjt/44b2TZwMGHhsEOS9yL659ps1
2M5KjgXTXkACKPXaQEg8WEfzSqB+6SLOgc2V4RWhBVsn6xc32Zz3hQgKA+dVTzRSOqZX+9qX9GD7
cRPlLzZ7gPfxQMgew/qrkxEUywvhSHULFeHt1A==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
t/p5VtZHjsLfCchUCgNeOz5ortjEuL5DM4rb5ngmRXsGy7TlWNvvGi7beiAnIwd5zTE3ry+PuJDU
SZYf1w6dgIZo6FrEdTzcaDzMVk3C+gqcEn6QDd0Ifwuenk87/cQHamfW/hpxeftli1PrbOgCMGQ5
eZPwaz6b30C4Zq8SPk4=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
geToAE9Tyr82BrB2vCZOkZnkALmXkgXTx2lBaNZqm+awCeqsPpqJRsQhbxGO5M1rnq3+Enuo3Ec5
RlDRcCjJvvQRicumzuJXJPDvjDiTDSU8tv4H1M2jUT5JIiq8eGbAfRhJDxmW+m/YEMo/wcRrzuqx
vIsEDAoFQl+5fFBytl7q2yYbnNdkwsyOo4IY118wbRAOBUYPRzTyLkYWkOMCnlF10iilmlpMnweV
wwRZRLWAvZ9TrXKXdb8QqhZ6PNINY5b99pi0gwFEKTGF5JwLigHSa41gHQEdecwwJS71Z/l9wew+
Lh5dkPFSfRaFyhaR+wLO+xc5H/ChiEiXK3gHmA==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14432)
`pragma protect data_block
UZ8+K5OtNt4Z2YW8Z6gFKR6IjRanOosRb6AP+SiPzyu0NoTuNPzPh5jzJ7Uan1u/gc74ZUvNclOZ
MS0PfH9jZOsDUY0svapeJsvSETw0bXZn5dyHlBjnmE4zrcELuRo3EFWq0cVkpkQWfd7a22M0+8nG
X8e/qDv5K0VM7BPIYBaF99hTxKRmaWRtyIuvxxLvnNY6WJ3tGro6dFecu2jTAV/xk0HnCkFyv9rf
2+wEee8EjEuI41G9y0kMxQWozxPQUIYYUINQpo0x11IOUdh0XVTHCzha6FX52ifM6IrUwkO/uODG
Yh/dqXWpu9ajsF7OgYRJU5268pFyExQYyC+pk0A0Zhf+mym25Etdug0gxhQOgX+6R9IqEiTfExp3
SpLycHEzHD/EK+fmKWropHQH9eBbBKSu1u9Zi2wryc0CZW3d05oN8TrCNWtDDYKey6Ow6xRP6vGA
DeEw6h4VMn2wjvXeYMoySS6E6cMgvjRcIjgJST3EThPjGaYyDOm5L1ChJQG9Aye5f7XAowLU7I3t
2atFL+mJAthCvWH8WjVbwuMHNd76IW7gJCA4yQRXyf+DTmCp6JSTIf08mgQZVwHuoDDM/zR03h62
TMiv8r6ZoSCL6Eqdnvm58tNDL/NDmjJT21Y2RrC9FLN29bbH4u0XXJZ9+A3juWeq0OJoTTUTye6T
cyRWOF6igeZKxgHf8ImMBC13O6/932+AKDtrVPZXq1fWmLwdso+EtCaBqJ0Sav0q52JLChamDC+y
pHuvBi5SmLJtNvL/ejB6AKA3FjQhPXjr74wRK4ZGnMj/BJj7rRiuognI+mFJva+np/DxYOA1lgJD
jYYJhz8ipCEqdPdQJw9Xz0CwTKUIWRk9w1OiZJlg+cfdAtZ757BjsFWun4U6v8i875caKV2IzK0U
T8zWDf+Cf9GijGNEYZULqjZhUZc1eGqBWx3xD09Z0ZVwQ19GaZQ0TrDsDv50Z8wKNCwQWgUdNalC
xugubqnRSLGXZUBzGqq9dlFdiR1ot/cQG3qhr1oWLMw4o64TlYBWJ9oyt3Zfd4909CBuF4uf8qqA
Ou+yhnbtQxujUZyaZwKbH5QPSC4bv2Pdg4MP7HbTuifoBPPqY1QCgtYI7P3JbNly5SIeLAXVLPnS
tt6CR6J3wwY2yFT7SVK3hvDMEGs7b7qEZQ7QqE2M9ZT+uu75ao9XO0uP5/p8lbjTZcwp2BD1NlA6
r68APcr1kw1lGhqXfYYbwRoEYuJ64siO1b3CjsLwHA4hlBywxbavRGg69NrefXIXtgNSJmPwJzz1
/eTkhicJWuy2y90WCxZXe2bW32T2ERJ9idqE2y61Df6DjYdyt8eendR2+z/CwM94kSu82t2+tguU
6UVLFIoDgnbvegyWiZv6j6U62L/fjcByXWfrBO4zgE2TxNc1t66zqDhsSR4yOJp43PqixHb0rFOq
iH7TOq80YXExLvjAibQr1JMpOmhraE6DGVxx9Kb03mjifTnTboC5ppwu12++mDR+winxbJ6jifI1
AuHcI1b4Dpl8JM71fnWoCuN2RR3UM8NE1zAYM21Bt25QBD7bPI05IQ8yXoORoOxePrv6+pROAzXk
102cyX2wLGmXmEOWADxVr3nTnpQMnjBJz9ODKWOENQD+ynepUUZ9/CSNcdpYCBbQBwfoPRRc0R/z
51/p5eYSsubhl3aSyySDPi3C6a7wjRdIsSDbiJqKaCqdt2bEN0cHggbvCRtC5GUAgjMdI4ffns3K
IjoznvtrfPssY+SOFiyG8EcxSFQfyxlm0xGjq75FMpjd57HzdLasM47dYTA5MrLTozx3XpkY0RrH
/DYxmjEFJMuCxkS+nUsjZBp2fP9Bas21H3BRSzSlYa1vQWEatIjmm3O1mG1i8iOHBb1sG9IJAMem
LAEbDqC1DHSWmcrLigB0wxU1cAb4RWSZ8Cr+BtLSfQ3UA4o+r8hU9XhNAEcK0FGss2hjtmHFWKV6
UcXSjyMXtDUZPh2ZgL/qNjbqbGX5/U0zXH70uPqY5e1vFSqjBAScCI8OxcOv5qhwzkFS5WPmv570
3AIQRhXAchCsWZg0s1mbmY8fEzrsA3RCJVYrT5/hT2uqgLsx63NIirS3i9REWqGzxm/GHEhZnqEn
zMKuC6HOtgwaE2nPqyxAZwLEXajAOaeWQXm/BnYFA6mvja9g5bx7fw3XCTM4TEtiAzwEekr5fwsE
uoVTpgzI5C7MZ3WAHlsbVfKZJkDjt7tCbVk/T0n/eNQpjjwB0wdniVC5D9NThsDU8/fYVDCZeFpt
MnrD/GAUnGw+aAUli+tmdBTjd5ys0vLV4nIUyL4L89HFzrSKhXDN7fr+08gC9lwa827c1yBpZxFM
v84X5c6FS7aiM2L88qI2bzlgu0scM6byBilaMa6u1sbEL4NFgjNHOr510RuX01Ak2d8DB+rJDyBe
oekfkbZn8+BB/ytbB3hLThSKsyPY3f74AbuvORls47Q6yAyjd76P/kTmRsJ0fIV4DD43/8xHKSmX
aZKoYV9gMNWGhIAF0ODfVPbSYuEfs0Awx8/MHV0/MsO40iqn4zxcl21JUgjESYIaZWWsG5jfTXlf
hcimRhtHL8VRoiYBd9VQEH9rOVXHUEAUKye0W8ycK1Ij3HysJTm7rPtwkCknhhQ+IqrDXNzOMe5t
zWbGgevND4C0Xbm5qsCI93Mk4d0n/lcOHmzzgRf5Mwvwgwwy10E6pOvQ+yiZJMdngKXF0qhDcS/v
Om5fq6JXjMt+voK7Kg2Bl6hS2g2wHj/c5eISENiS/fxLiYC7JcCADUK7mWzhrOxRYVXwLGGlWvOk
84wPT52IzJOWM7GDbUSnG6GhizQNrfUcf+2A9eM6bqOmLoP8FL8j9+6yD3JIByeHn5YgSHf2zSmc
RRIPZvhysKJ9uyeSMb6LZy7QNbNAR9NqoxiiR28uGJ20QrSSvU8B45urOeKzrANUYBF6LnwAQGek
8YC4g4yxWI/YlO4zhn6dZxNHS+8rrPoCRke7VRHFOTD+96iQ0sn0AhYgCn5m/QBg+t2ayL78bs7p
kx6s1SyCZiPsRwdHLkLyXEk8XBP5ZGhYMpAcEsBGUKj/ZJxuxaweIhQzh9nhcFGeceVqLaX3BJLp
73BGVIi4OukG5ZJ/qAjU3WwjHc8gDCAvgm6dEDfZdhcFH6GZGC7eEkbuyuc3A/qD3rdqOkn7fTDj
F3UT+FyYWtRFB3tLVxkSfSQ/x7SxEb6RHUNYsDzYh2K6Mbu8FWcuhmqT6k0hxBaULoRL18WGdaki
8uL/X2g9LS3NdrM17wxZ/li8DpAAUb3M6WwFTz0BdSbmza/Oubk5XY0RLVjjCWncSqihpeI/xKLH
vBySDxjeNhSrP7OxLOoJ0FSCNK8941aVYOHIXb/IJBsX62w6Cd9lKy/4TJFRjihdjhMbRuzLVI18
KP7p0Ja/beYffVgQ7mPORJBsDudAJs4t5ofl+V90jLUh8/9oDL+hH36qE6VxNsdYitoLo9TlAA5/
pGQNG/XjKtW5X9D+DwL7uBu3F0E3etY7tRxIPjf81fl3n5FMZm4WhRmCCut3F95+37c4ZDn914Ry
pTPaGBpjexjpgOKRPL4EaWZXE/IMQ8DBTBqDD4+4cBpku31nRZ2KvDu35WLQDYfTaC0G3mMOoAEG
SKTWmgRe/X8qLxXIHZve7cmfcNVTAk/J61WTx4FrR2D3vmZPdMTOasdSo8/9f+NUyJkyrNXO85Ci
1JyVpXkIUftrMUmsAePDtnrsktVy9GLjVSU9cWDXLFde5COZpr+/TtuNYZzZdzkFiumV9FpKvgId
y6fsbnac2ShL5Qr4N4DISDFlAYiZG03kjcnsWUrtCvLNCThD2zwF8gPimmopPulTlLt0KE2ajBsu
sn80gODBM60IE4MBTJpa3Wwp+TOqPAZ8iQi5YEaM5cLjqZOTHAujQIhh+KaOheODnt0uZQ+RtFTx
829jR+is97NYnDgvcUVq2kjKJ6PRHA15bDD0UetYfFlfa6wrY08SQZ7gBtMOUJVv84Q4PP+uDO9v
UkFDZyyiNiuvQEec8p7TPs839+b50k1WOq6g2VVdRiAoINuARPQI87BRjZDEgD0DCgRjTuR7Vgz1
+yBojQEHbLRMPDEizzdQlgl8R0njrsmyFkVQhgUbZDcfMbTUBjYeQ/kY/zrhbscYQu9hJGXwoaSD
qUuizCNQCejQcUqEM9MgTAwovOh0Vunknf06wHhCoJVYkp9m9U9lZS9vY7ins1DPmp/Y91dOqMOR
PzIYzI8vTKQgQ8q4WpPgKKLSZsvCUS1arUWabovr/uhDpInqTrRPDiNSElShIJdB5wEd4waG2vlF
kKa8PsZWNAR5c3giOvoiap2UVdal5AWPjBVvttQoq+aeAOy7bK9LK+Q0gnKJeuG9UGbtV93CAMP0
8vwixyD0tN/Gaj9p0BtLLKTeyie3iniOUzt+Fgd1ED1tzQXReGwRGYLlBajFid4lzJF3P/VE10eP
VBJX3XbRz82X/ZqJPYy4Ifma7YKoB1GJGITtHO1hD6ULtIje6G/EpQyXa5/WqLDd9m9ZegtNKaPB
DSy9x5r2IJm0erMrYCcE3FL1RFeTAolUQj931uOH9fjZEJZx7zxpA2ss0s1kfUopAz+7xhRN0CfF
G8J0jP2ZXBS++yUsDnJBoBBY90QglHCo5ro1VySITKuN/1fpjlsFrACIAAteDsbsKpHRe7bxEtJ2
3CPYgiBq8DQy/t6CUuFqHZ/iR+AtvFoofR0+GSUHHoKHfNMeqASmAgPSwu1cRZYnJGmF56wnwJ/p
87W+reTMaPfw4dRQ1nh/i1dMeccOAIahC0bLe49qdzJl1SAjsU2o6bTo99AVl+RGWMotnYwsWSxW
pB7vR2ULztAqmA+TjEbimCZJhqIEeMnLyI8iZLkdXtXwgqWL+1IppdMP4gcrzUCdZ9XwqA/Ze6zd
p4KJyhxF5O5YYuLk/zNF5vKSfKSsgUWF2pwECi1j5ZLIKH5q8tfb2o+INatZnADu1q1TDfuXR0hp
+xh5P/ZSLZ9dysGYpijX6n4x8k26SwbAPFFqLXQ2NpW4uMjfDLi7vKUwt+aCA36hyHNkHJfGzcRE
RZW9lTMouyo6apJGyEiS9qDQUL9rJcQY6cSO3AVtSb/a1h2Urr/GrkgBnpv7HMWkZU2EMwWfNr1G
jAkIgw31zrqZxHU/UGr3Hbf84JGQUiE09KLUff/Gb8fTvpxybDsNWvE23tZws8eRPXW8miOoGJA9
xZQrNnwnMZlMK+d+m/dtLwEEPvX20cGfomm7Ws8D3adIP5sVrZe/KpxU2kv8NmHe/dfgalYbOYfs
ZHQTRjjg6URuqbej1zHuH53ISXeWmngrIMUX8Kx4YYSB84J7zYpR5jfyqGTIYkVLEijvbmo4iVC0
ovdWhhssBcWOKvRSjrSiOC50wTkDkDk5yoKZwl9QarzojxDt/t/U3wtcJq+cd6Bj03mB+zVPT/0J
W0zw9yM/vWVk+fIFMXcQDKVfMi8AcHOkLoFrpfWzbMpjbyknDstdF1lKTwHNRORJFLrMOQyrs8iK
xfoevI7MQ/rvoCMggeXgswF0x9ngCCbbrdGmeTMhvSk5dEhYhQ+K6Gq34ANhgZvBv4SN/AAPTfwH
4mk2SWMhCqxuEvOz7gc22kjs7nYBAhQaXL/otSOM2x+KGUu093t3E79MN2vdZqXZbcBSnxzM8/F5
NzTRT+OcpWgpcaN4qEAMKSHedhdzlVMXHv0aDMZ1p80zbRDTIbPKfxUWTpq19ew633gfoYPX1SCa
SnT96VJ1kIsKRHeXbchZAHJSybiUyR2PHxRPlpWpww3321g4DFBCLrGn3s8bbUdQjBejznTThsvo
ATAs5q6Ek6dqcwxK4pBUXorIajAEQ8asuWmmAocmZ50nlJbsxfcBlcSSKpOMn+rWPmAQa+tXPyzr
vla8YiPR9HhCg2t05l0wA1+3jFEy90nnmfCRyQB1K4wUN5tiMo48C0QW0ihVa41SeILN36mKBtN4
TNQYke4SKb4NwCX6jRR21fybXVavx1cPH+NAgcNl518Ir53WMmPfNCz78d4elEcjq95q3wnxN00V
MrRMlzneNhWycU3ODFWeR0BDUwo/DKEnEcgxiPpNMHO9PrKZIMKG+dVIZ/DiloFggbnX/3gLZAyJ
R4tDH0xGQ9tZf1z8G7dAIjBy/N9J9/iY3K12vS+27s0v0BOF/BqmRs1RdVAG+nYjwWJ5QZokEyDl
rL9ie6RXq9Ac36XwmYFzj/0Y6UItWCCqH5Y7Sgr47viaDaqDpNwcffRjEcy1VJkFUiUK7M0TijT6
rYvL+eQbja+aJY0vZCuaGrNmxKEm5O3er4PUXTAZK3T+6YMdDUh+qMREhPAQMGrJhWM3uibNBtz5
PFBSoBpBxZ8NQjLdbb+wDbX1Iw040PVKJ9D138nVerpTI9uBhiMuyht1hWhVuUBNhZa9RdmAx/AJ
BcplwYs934hkIp81b0opgeE42wKKLvtZ5zotvNYea971D9eOSblDaOQdlFAdptmJONrvcww19Yyt
cC3KiNeBnxI2K/CJ5wuSqm+diJZbRiCH8J46IgGpHMrKC5JymLB+AazZDhmRhtAHJ+N+WXbBpeAD
UG6jcolrytBQJKBcw6FmAHhpUQduZ6pshmWAztdHCLSBYhziRfOrt/hVBP7Urq4ith0wc6U2PpKL
yVpWlyvhiJb7+p8Nr73xYu47dSBs5BY3hi/w5JAxSMYY6rgcnPEz7il4V10Qc/O0lOEJdpABTxnV
iZcSogPEZH2pZYzeTPWlb4DJM+x8iNBj1e7FKVGrgJqakNgilokugcJWMjEj5oGludiiMuktuRTp
UjlQN9lPWFsf+6zWPmfDj4iEuoiTLqiTESby6zmKc5FQnfnpDEw3bb/aN/0DQ8Jkrbxe0R48yoEX
tt432HZhnPjKQiCxDYJA/EHCW0Zstye3ldc/7vJuTTcQin4l8szMge2G105+M+5vCqQ7K+leXBTZ
2vBFmYF9S5oWGvaLs7sL06JDTyq1TXIv0AMz0Rb76lzxQwHwtNF4qPn8nzMsdPgw6hl9BUE6a1mX
ZmhShZYBVGEPlA+DrPU0dKliYMofcLpF61wnuaHNaKjHYq++upe65fMVjfI5kHPCM3EMMON0s5Iu
kUW3Uhm8f/TEHiii0aNVZ8BsXcigz3L1jdwnjz4uPvH+aLAIYxeAv9Og5zaYtb8GKaLeQJ70IMq5
wZVT+pczO2StE8A4acWTo6ajGL9soI4kXAheog2prnJGJi6A5cwoDORSh5sSbVLtdcZWt09hzWWt
tPemb89MfvSzkXMAWk4buXUH/F/YCexI1kunqbrn/U9ixUiD+HtyyoY6Tk9Ivex+QpWo5je2HJcG
MW1ajS4ygOWkZscenJ7rd6WJm8vneQdGRX5H2oWw0YmCbitCY+4prqYcLTnqt5uLbQvNovqBHW33
O0msV7Mebx5mNo0ey2q3+a5AdkoIHP2UGQD4Np9IocPnluWd98QjN7ITdtqwCsjA8NgnHgVeg5fw
iQDdBRBMKjFIe2V/mWol7dyEFd0EEYCq+LBia22cKCrGPeLCy14Dy6PLo0Lw/1YMo+qPD6CcvGEe
IdOMmC3IEE2/HVKxMv5VRjgL+Ex7qFXgOCH4v0/Cpb1M+kUb/Bz9JLfxUYRAuUtYqYvrnA9xNT5J
wxpj/wOiMowoxAl74kZshcUs56NHlKcjTh64TxsIzCScLrI2LKyL9xyRSQ8EGnTeOfrEZxucd+44
0alF63/cDIWNKHt4mOYQSeetbuJTnC/K91U/TVH4cjKE2BKs7syMo9HT5yKkWVnsnKl098Kxc8W4
zvE6HjQTIxY0cr0rAIiDiOTYa4R7/kFj24z0HOtNGOkt+NaCmGwo0Agq4Wka1BNbK+nKmY57Mtcl
CSMb+btnYHiL9+7gAshzNDmqt2SoS6kYNqzD7VKYIxxqIMIrSCr1lxk1fxpch2IzSTZiZtjt/hTX
rlyPjUvOufQs+ylXw2CD0ynGJnwsg/fnN9FgjfOLNlKTvaI9DVfgX1Qi7RjUjO4nT7McJ9ebekJg
uNfVXlwmnqitGhbrwqHA+VqkXa1afFrg+1VvMKHoHWLFOoTnwZxAsjNMi1YFkk8qRUVCD7FOpEMk
Xn6xZbOvRydDNl+EBqEXvX51AT5N9TTFDp932YnAP+eWRPfqx6GZuMY36VjLcdq+w7eutcoVxT5S
cTS2F1+YwEq3RFXxZlPYBQBl9e0A90J8ikSRKHGF+LdMpUwtE1oGhQrD9pyvDsPw5UPURH6He3BS
jjFT5DZo5YIhcZ7Qpr3QyiEPsSy66/P6vD7iMxlgeVlUG/iRiOSKyqWJXd36ZN1Xjum/6tP8/Yfm
6dXO+FLZF4LUW8eCWaIlX7aifdnH33PqpwdFAjE4kEC/cvf5hZgayUEH5DhzgITr21N9+20fR/dQ
R68cWPE19SkdC+iGuxRWW+mfoZhfYoLIinJZ11ShDWUdfxCM5yZ7aze7/NUlydDg9cfcUaIc7512
3QaCIFJtqGVvYcYUspLhQAevdkZhnRvok9CIQ6KINzsFHVKFqVrNclSif/HfspAof7gZ464vAQ9U
JulFwbEGTc8FpIJfy093f2dTcQgDPMuAZbQZyaJpasWYQvS/mNUoZ1hrle9O0uh5LnMJuKV3KxXh
VpUJG3rBGtNLBjhfnE4GKv0GLdEh0xG7DxS1AlM5XrTW1muaePDEyEDosyxlJOcajQLb9OyFdYvF
FN/JzhKaUDCo9TugUrtHltDVr0iVFYwBlFHsHDxZb/BHHe35IMRSfT8jjDw5Q6526C/IXFaXW/VX
bvZsX5m0QTf5yxbKIahBlVUbMRpqcxClkLsqKY7fWsnBFBCSTv/ZtVDARhEiYYO82QQacH1i8RPo
uE0aCXWspn8Dp1IJ0qjMG8KdHaRVBsZdeBfkhEkPdyMV8G9Yu0U+rJO6zE4sv87YZvuyMT9fSX0u
WquHyuVpofc4jHk3TQ/1DCbtDtkf8jq0Sd7ZubzMoS9882GoEOtKP9DGRJxHlh8qIglNLCxxGugY
bZNlipa8WZ3LilE2C2SYGcJIQmr6Lm/crDVjAbcnuxgRYJyhVz26JEq0/J/zT6tQuf7EdkBQyTRe
xJ9J0QSLIENywec8ttgIlgINWoyV9ZBwassOorj67kNuvzbs877gbs2y6eQi0Zggu7RPSGtFG+Xr
vrdbwt0+xTWeF4SPliQuKtvVgaWO0s5k/KJ5sUlgrAzH1VsE/R3rHxM0QKN82J/CrCNSY1Uugqaz
xtbNSNtSwgVV27VF8g+mNS/EFxFGPM38yPL+dl0yZbgNRiBiXasx370P7/AIAJWbDOutWaX28GD7
W9L+TXWtxbK7/c6GqK1FjTGOZWVzbeShcNEknCEVvbSIkGrlkOojnJEYzGBHH3C+M9wMb1PXQNxD
mrVCSy2G0oJPTKEOro/ZWqq1GyQBb11BR3tBbb4OXaTXKgZkaPocKIdUxoIvqTfWNLszE+xrkjyh
bibLZWYUGA5fcqTE3KmOAYIGo4/129SX+FOesEqq8QxOPK0c6sUv8TeJM/45yiNbDYkNRcJe1YkP
s6evLVsxoeLtO1s0kV55oPUQU0CDtBCRn1Q0sLZ/7S5tcV5Jwp3+67qgQ7uFrzK8FpW30igPWj71
UT0zMrtQ+iAm5I6uDievOTOlr8dmPprXyUp6hRt+PakvQxtz5byaNNi5t7kBFxXiJ79ZpxkbjCJ7
EhEURPAUlyMdqD3y5VpQ9EZoN0ftlxzziUDk4Dghw6PYIojStI9BNNIkIBIX9P6zPCfBADHnCVkw
6HdKpU7MnydP7v9XOsJ3Y1YKUC6ltAGnHBadlLQzsQK6/pM5ZuQ4T0n9b7/bOcwjj/I5R6qQ5Qzn
PWehnY9sexfctLCecUB43P8IWXulk2PWnsImnzP/5wYFYAlzqsj+W2EvJL5bqudy6JBsHOjEoEll
2Lcp/hyt+ZhTPTbbsmZCvrBp2qBz8vbFtvxUbhkAhy2hQ3qgX3F4J+m/4wjVRtPnelm831edb5Nu
GrWHam6SL6lyiAa+CNP0smmc9oAcvNSzUWGhbqdENRtz40nPIneLqzAaZj0BCXFzMmdCINFETMUn
grdWC2UCXWh/Nogm3FLqu7+5US2CgR5XtBRS5tADaYuM2F4hab0jtRp08z6BDUDgBasP34BMRtmY
INZx/7ixw6vLM6myLkILfNcPq2N+2qeMAdjfj3HAKQK3rI5DSV3Rx5y0taeeaNlkGpb9j2Jh0q0Y
hXUu+IYlgcf3K/W5c9vhpkwXzNb91tvgVsICVsRzi7Yr/Px8wA6fmy/ReR4rVm85+BjhGmIOnFXG
i+Bs9N6LJ/gnPE/u72oyc4/igWEfshrBgR8+Tt+FAF01lJxmbYvlQnqFthxXX5TkvTQRlSPU7w0Z
u3lm2kk1Uhx5C35EnnP3zPdYjrlBpGpz0tWuwXaW3NHgO8P1j7UgZJAu63J6Oz1VApYdMw3TqwVw
ZrxpT6sZx8kcF4q46fiQXuw8XH20ouxMToBrRjjYTrlZjyA7gK0eEr/+BVQKUihKidfUSz4p5wIR
PUafoOABgNhE/igOkNZsmIAXxt/ZmOthQdo+mBoVBC5uHMj8oBYa29xCqN8AMGNxKN3ps/+LPUPg
odX2wNTvMv/JebZEy1cnCeFoEqSJOwymevEM5NIE31f653FQaxJJ0b/qXx/EBTMDOZZjqI8Ahpvd
0EoE3SfHCDhxSxKnxLiktUHwmrj/tNzoAQQfPsiqoEUgyVMGP9IFC8qf2NKpqsb8Ov/XMqrUBrtL
+JenuzZmgSJ8QO91YGashDJtJhC6qHPMCwBO5rs+cjZ0hrM4bp7DbyICtHnG140UUloROQPYNViS
fzmC4wlYzE6EQh6x2Set+yQLaT9ESTXej/IUvWXrSc3omHhEpnwlIP8m5VdKXc8rWqujjBZQOyR0
gGuFoA8U8/9CnZwn1q974k0YwH0CET4mKDmhh/FX/pzO/YcVM+gPEXML/F7qc3Qw3IFREwyyi8FK
K/i03PtgpzCS7TufduZXWmIrbgci6wd0rZ+KKwIHMTUPdKoOU2uDoIgzfAAD+ejeUzXCQercu8ut
2HIGNT21G5faFrRu/yH1B6iQA0aU6MRmE1uzSEUptdSVkVjE5Rlhls9aVZIrkJWXnP+ZE75wbKHs
fbaDoGEKVSb1x1caThJRzaf7hLj1KVFNE+hCuRBUSb2JPle790is+KrWbdfcL+mYZyPeWqpNriSS
+E+3VlG2WM9O3UP3wXuxwazEBP3ldIYQWmVaOGU11gK5Hs5YgOrF56ZwNCizEyiRrGPh4YCvWr1N
QinPrV4EGFu1lC9AGYQrdKGHEAIV9lcin4VaBkdQMXcvjpNtdOcZ2dZKy2+Y0OeE8aI2Nq1WcJv4
ODqf3bmCa7WbkSg6zr4lmTIgdVoUxqlKS4bMnccHZ8UP0P7itMf451M4ondanJAFhQhqQru+xJ49
gH89VG5ooURLQmZC39+IHZtn5+P+SY8B22DpTvmlALMGqcLniBE4MkLEhP0v4lXnAMRm4L5XbChz
R48VwZbjXf4fyFsAWSIU43WZAGlxsXjKaSSuNlNH+gta5DNp1QD0gnx8hoEgIKpmn/bY51n8M49z
fnbx0voQ+R1CxKN+H12NIveNkkwNscupyuiLOqyw6vA498iBFHGrVvR4mE3J6WnLhot7SNONqivS
ZMip9Jb+hBeJ8E5WnEIlP27AHG3TeE5MI7IP2nc2lV8/bWX/p9nVPT7407ZwI7FTNUy8LprPui4u
iJKaFMVLmQcx/DbTOiZchZl5z/K7wXUz5HM2bw+cdx9SZlHILcINS2JlCwpC+Cfm2IC9fGOGjpVT
rgvf0i6HUPUvijC3lp+cjlRFXdL06PvVnvN3+I74Nem4Ox+Qd+odeb+BzupCD9uWi5MHSx17zR0t
yy6Ywppt9Ri+y2DPyAB6Y3K9gG1Yf4fi+Rbiv7juCtap3dm0ab3I9t+Q6ykKiADnvCvAbdFmWL6R
166yUDCgTi3mJ8hdj1/0ljKWFYWgV66QxY2gqAoynkQw+Uy8l17tPlxDSFQ/R1By8pfOsjOSEsoZ
Yb+sf5Hb1O1KtC+C3sNo9dDk2xIZKy2LHQRQTwxO314SlKecbQUv4IgOHsh9oj/7sBzWjdRJmyGO
ykNu+o1rcipZPBT+EMMdNjnZUEYsEGwve8OS5AHuKVKzVDv8CV6e47KzI2I2n4qsLXQ3KejPRoy6
3F+oXoCYbn39KntX/1SP5C5Tm3ofXxh4sO+G9DViEyVA4C7u5edyYqG70NgfGip84l4yiDu/BIXp
svoZMwIzFPuzpKhEH1qOx7hVREfJlkZneuI2mp4vz9F9qGOOGS2XHOdY+eiOE6UtwjRyn8XfvTbD
BS2GXGpH5SW2qnBZPxTuW7QmsPdIvGZciN9IyhKgtUnHfz7FrhrDKtp8v4qpmlaZ1VBJd6RRio1M
PA27rMAjWW2QoJbk29LUsMpoOZK9JrPD1lYuL9y6TK1OMcLDmX8jpxjoQ9hfZObVFvn5Z3E9Bply
3Sd4SLvfwJmDcZglLgYOCAuwUZ9YA2lt0fyvN0Rj1L5PDmSLxr0HFXi63Y8UHPULLctj1g3i07S+
oxx7E6di2eDi61XnKki0oHEWH0ork0HPwv/qYqQK1VTx1h11+qV2WQxtqRHQieujEE4nPtt/xxF+
HA+xU0MNl9xZzDTVEwRDcM2u6nqlZTZmJHtZHvFVofxNiKKVX53864orb9uIx0yM5K+c99h81PPT
a/qml86+xIEXji8o3p7V9xRcIEzigY7SeR822M9Q9n0JRswi4otcnOJ9gHiU3GihWCsOwcr5nqqR
gdpYluLNUn7ZOOhgXaN6O06ksEIVIWzkGoro/GcA5e90sltF+U2m7XkJyBj2PJ4JgeJtD2AeyNrr
vXTiJHuFXtJfmDXJdWVa0gZIOZcG1c+0MzvVBnrCj2ootAsCpoVncRRUrIKE1GwMR9tSbZoB8Nxa
yG3pyeimlyIJhw2EFq8d/9eLrm+gE6gR4AUW3tqRQV4K7qsC3AJ9dn0Hw927tZ2lbED99Hji9g13
GcMUroy+hvi/bglvl6oWB/vu61/a/v/UEwrCYKGQequeF4ts9T2BBmK49UnP0NuFqViUN+Pqesyq
ap70NKZaQhlE+tDNsTkhGT+Aa68HsxvxTno1IqmtLMNno/sGHOb/ntT0WXvlj/GiLMWXaUXUFz7h
4j8d6gQn68SRk9thR8nzgDA8DChf/qxe1h5JTGOgyFzzUlvy/pgZH1CmPb5qa9UhjiJkvC2DeoE3
lTu/4NbD0dCLia+lKz6p6zRw4WGo4PJ/Gxg7ga4064JRW9t0zEtLKgLssX+6uDU0SxouH8v0WyFY
6TQoZf0Om5xQaZ3iUT1A7MQUBC35ywo7zLbE+U0KgjfbD6bLxN7Vyv0AKFMi5m5HeJsfpnVNe2mj
gDAY54dNJS0ck3kIHfYExVtHXgw9Jw3IdntnubD7WnFQzvANkbVWL6C8tB5w0IDesi4/U5I0d7DB
WRPU4CQMySY91JUUQj/BvL1D+kWiGtX72NkzFq41AasOwc0XQgk+aTIGiBIX5lAqNf0BRxcPmScy
BpbqIUjQNggL6K1l5YAdE/bEyK8Hah9UHjd1injRrQDf57/vZYAGaWtYpI3JZ62LXDAAVkxP7Ojn
Qr/F/EyL2cMszWca2DfzTFKxOQ7ZsNDqQw3rfZhHnXVEn5WJVuZjFkRb7h9IBD5Tio5HZHhDjyGD
Z2P45gDaMt+tNjn4J7w836RCOOekm1+63448hwZLSuUm95VwH1BlaYwmRMCIPQyAeBIz9BLdf82Y
VgrtnKdjVcH7d40HSTRiFd/tFPyMjfF/xhm7boq0VdOulQDmBQ8NYKUhmgY82iwqaDyBmL2a5qYi
mMBoz6aQ8LV4fwPP8UehaNAtxQnlCEbF77uw4hDQpud1oTTFKKVy1tINKT45sTSnqBSj4WRDSYQk
qtuzEQPZNwH1dPANTp/5MxtmzHxqyMrSpShM1xP0qdX9HrkcMoxJmRT+4JoMI4AjJja2+3oOLUx4
KVBQh0n9jZmilsupwodTy2YW9snB8xT7reQ4XzhfCUyDuQSm5EpAnJK1eMK33+KdofHi6qmwjvbO
bHRNWqRuPSvF3Ow/Nu8T+A7RTN6EMOmkKhio3q5Q0GYWUL8dFX5ixcPhuQ5CDFLQuvsA+ErVfWwN
hO4RDuIe0vXyDkqw0N/9Xp11Dla06gWTDq65YBFUXBt2q+cBFQUqzCeGbI4I4ZMWlvmBEm+G3DYg
MnVf6Sq7K8Q619bNYczQlM1qVsldaiJO7u1QfLgqlXjiBp34dU5Dht3ZGrusw3M16/PB/V17uhf7
rKGlUZML0bolI3majt5BTez9C/KLjDoORbJsCiZyhlMPvr2F7ea3WlT/TdRrijlI9S5FMOBo1VzQ
9nwXRQRZfy0t9efT1RTcpJblcl0QU69AgODwa4oUDPzityZoNPPgj/WMgXkYVU4az5xE7rQp5veP
pXtPhIT+KHYzR9GVmE+z4fvho4Ekxwg73ivXTu3z6ZtaruKz6WtNnV2snceFqwLk9QZnXie+4Htr
gGYWIqePOsfQ8HKndXydg5jchfKuCTk1ugsYPaYXiVlZvI3vvmB+zSYDl/QU5NynxWqUG5A/Q29h
f+OJhXLHSvl/DU2YwhQ9gAW4+boGWj4GaM+ULk1nwt0tpNbDctsCm1FgY00uocT/Fm55dS6UTe4y
1HRergJa/O470lSgdtIxi+mY0PfWHNWEjJ+9d3Rs2BhAsGRQOh7ik4pmAWyZpkgnjSFFrlAdOhoS
CP3FXEAGdsx7qYe/me7Zl7JoKB+k4T1YjJHrGmyarDO5BoXbUqucMbxlHFZZpLu2oRXGOrTX0h+7
P/o4MUoNl+7/btGVGNynxbmxgGymflLkeLtV3rmVGnUQs/iYhFYcLyw6GKG6MzZ1w5UxQJQmYBvH
/Yubdl6jjwXGQEAHh7/62WUzhrpf3E8K2Gb3ueXbR5jMOwaO0LlIHmHioJEsE0VuIhOZyBx3dAau
VHfGJIGexWByuDHmosvEYbKJJQTzuAuHaNXi2fXfwewioyVcdC5Z8GcuqMCblD9b7r7U/jfFH7rd
w4bVbLCdcVd1HuAcnmVtpg5fhcTsaIZfd0qwuHy2ZssToL4V59Kvys5GPmxcKOXZm0Umt+9jnSV5
cZR55hwUx4XgbBmmNNzv0dE4I+lU/unpE3tK7As86eFAziC4TYNHlYfgG7D/EaUyYKX1agIZ1pNA
DOKbEj4Id4f6fm/zDXUedctUuN1sLluLq4voNM83S9lUjgkvPL+DyUQhGCoCbeVXAX5c3fmacQw6
GvBticCDOd0FX/AJ4UwacEVCWnglety2o2XTGEZjvT0PDsuxO5zZ7XFjoNrSPj7IUEdKyCXaOs67
qHTu0nSpOMoRyO7PqImJpTJew/vtGvb2/mBAJwV+gqhmdv0Cl8hSUHOSTTY6qkANNXflVMbGv3OY
kwcjRvAyLMjaxAvhYnT5gq2hCBNJGWfhYlFZWJDKlFKjkzb5IVz4jcEBCa1mi14zfZwDeciIy76b
VDgkdAdRVgNsQPGscPbpYLPDYvRWkU9mJKhZdrnK+FNukLI7GsQ88u0NFXTQKcjwfNmira+mu7ME
wnijMr+Te2D+4HjCnj7HMKlkPbEAT4Mp2tU52A2W57zAWeV+czujJqODMG+kDItjJ2v+LvYnMULg
w/bCY41BC9ejv77K/LJ7eElbkXU5QdEb1ywB91w/VIW0srNE0ZjcItX8SeCOTNIwUlCFr2qlg/ys
VVKRdHrlr1rX+4B97AK/WpD+SGtKHPySeOE9UIG06+6JkXH9WEHO45FBWr4HmoHcjXSrn0ulEzyp
ZBzyg/IUQ3u5WX+RbkDbFf6oWMjaFsXOepjcYHSZNoEe33ktqd7zTdfBqqnm1j+fY6+eCZSubC4W
IZhFw3KbIkQXWq3Eqh892nnqX72Jk8A1Lf67SVvtgftv+nnbatqk3//WjmXKRR0f39wycWCvxXOA
GF2VtKEYc87586BWP/0ysJf9ekkZy2OuKfeB/KysZo32L9GNnc0bsTNPFEymqoNYm8EFVz0u3otO
0bEpyn/qdJ+F8X77wJjLWS537gpoWclzULYWaAPlSKAO54g+W1hcxevE2iz/2EaBuFI8bRxSMp69
E0NGloUG+xNoI2ahMlC+nO1SGtmt7iXED/FTnjSh0Hf4civYomuMRwm4iRAZzab1A5ucTcI3efcN
+c5Km9Heo9E8WqLmj8UgCa46i+J0B9oKKC9y0q/R0vAt2Abg7Nvz5l6bGk5UyIAQwIv9uiuhTA4y
DUq3eFhiH4qVsxi9jmVeAbqUm0h3VDvpI8IEuPTP61CWgo3THC2syHIEP/ooYS48muEAiFjiSpvJ
VJUUWCtLozMf8EaqFDX1v3HxMzuuVi0NvGny5WfnYBuezvq/RQ7HxLdOWcmK8PRgwbcZRhG4u9ZX
I9hvIRcFu0aF0WfiTo+pbU3h/rh8GhJ2PUaprc/boqF+qWXHH+BYyGK8MARR0hsgs51ekKwByyQ+
FDVJ0Ry+uzWBVm72PhnbJp5yCyi4qP8bz//NYZmAAkf6KjEs73tIwFUzYfV+CtVALV1xUtSiMMjV
QpmyVtjs8qzIbOObj6kFG4iWkfoO66kjq1/KEzXj9DJ4g0pjQQ8459Uw+f0Pia/JEiSPUZFATxE5
mBzG/bGF5zpxJhM07WqT6DLOEUIpB0Cr9AORx0N8YYlcWS9kNGptcabgYBV6P6VExFb4spyNUGsD
W07Pi4vsnIn4s7pLitrwIYdTz/9vDM6HtF+jzcMGyFH80spp8Q28Y8Q6p+UI5NWX+T8yZaFwZzkL
GonUIU8VNHFU2OpbFJjRUHQmefy1JdwQFTd8+8qV9fQSKwo5hCk2QxpuKYyrWpxavMOO0wEwCOgn
dhtgoU4Xi/bHp/zgcIImg5YEVCYu+qXqhJX+798zdI7x6QMx4Jby+BGbc1Tet0YwFCNwuuArt+ZN
fN89o5sua3iWz3HAVb1mIdunHZdcRJvM//GflR6bxdzSmxghV+q78v6nO+VLObkCbzsy1tLeSD5/
5CADFB54ovQMUanHxMNVXRXTa+xeNX/eCc985gNyR7aN40nK7zIYMCNtZvknWXLB9rUg1p//ku0P
Gt+MQIJVgAJ6dViKQogHN/EBB6CRZlMXTNi9nF0sg84tob/HJt4Ro5fy6j3fpqZBU8H2x36jZEY0
EW5s/WSqAqFatSDEOOTdN8vhqCZqLIv/wJrYnfiYpUiYM2zA59wqB69v6jwfzsytf7epY1IWzUWO
3NM7WkCVrSQCv59RgXfK+6FWYygErllRC4pzUDOOzE4xAqAZh4YbnB7vxiqBm3vA64uTtTfTJiF/
SDkmncFHHwu84kRbrDQxX9AJ71SqV74RV7EnkuK6MEW3QQ3gGcKY4TXpkR08hXKCfR2hmgkPPd6W
9dTDf/porBJH3vzQFgg8GX5nbby87ztARUFxjYWgVRoXm2j+XFT45ONpib05ViLXBNOnNBCrFoaT
lOSQptRv5NsT0r5QdiRxcUdQUec/PqFYmhVij2AHUbD5oxAtsJmJZ8U7ElFAU2eVfsKQkiu4tyRS
m6kvvkWPO7mGnQ0E/AaXgFceOZJNtJbuMHj/URXLW3OIYnxj0VuFuJopl6r6G6D16NiP2aiz6qMn
2KKMZjUZrBChLSSzidZHfgxva54dTG3Kw1AjVG8vkus65L68dWgSdfMfxBpTvbMZwdJdjZ2zuHsQ
WQBPX2SHTwUiEmgSjH8ECthZ2i0GbgWGGVKcvUplzWtOSFhMekVOLIqOV+rtSdfwcp4/KtQJXxoC
FlX3RF9wZc3S14XrVxjvPHtgCfKz1F3jjWad8GK5rcw/BQyaeIjQKL22kX1gpvOn6NmnAFrx67Ew
7RMNlAx4FrKvR0hRUkrHGC5N1D3grZnRUEKV7ek2pUOLUPWnEDAjarwnNBHk8Mi10yLJxkrbnNFZ
hFoxANQcZpbVsl6qV1xZNq8R+EBEHzT6Hpa+4hQ+odvgxIqlg7szmI003T87lcd/NhlW6l/V8R5w
8bmmvrlOLuvIcvYbYHzUgyu8TYt1gTN+h3CEUBqoHTyOw5W4kMo+ZHa4nfdq2Y9730gmkzT21orA
S7KDZKuyhmlvrYt1E3fswma5ZATzp5348iaqRBta38d+AWW3s0n4fcgwtlglwliZ6LQalVUfw7pY
/3tGoOTczI1gAHoBei3Qy64CJB/Z2uZvn2PQy7MogsmYL0DgY5KCJiO3WyZCo0W3RJ9toP7LkxO1
eNoAB0mRv+j5P5MEmcfTbSaC4oHx9ZyDJzejLGWWkx9YNgfBNm5Z8ft0Szb3iOJewjfjkBa8QClD
HcIM2BIJJD19FAiTD6t/Ltb5+qv1UL9xFqfSayVUfKUAip53/PXHSh1XrctYNdOAA37EM88X4eBu
5KY9PyPQ5jRcLY0kEBLVC3k6j6s5qFfoqNRbqTdkQsKBrOOK7AcDMW2oW55B8zzVFLSujIv4IUpa
YlB5YjueNpgSaSm/vAjPaGTs5ZdeTioVwpikrb3sfgCqg7G1owCiLB3pEQASJes9oACp6J55yhkt
WIokvVqYEmhWIqs34cwxtVEnwkMs+IBo8Eerw9q38glkPIGE9WMxRiBb/DqENKHHmn1i64yW5EBP
MMJC148v7T1laGlFLcQGqHR8NshKNkg8Hjui7ewN1ed+F3rcD4m0qa+6H+rEGCuAh0VTLV568oY3
DTP8VFL8+Lj+QWUlJYG4Xoiud6KDWd/fTfwqsiLwpZOnv5iFopsGDbvTogw3hq0148UxIfW4X10M
oWbQB8aWD37S0Eb8ptf1NnE+B0hOIjvGvGSejHs1Voh20qy3BRdZmiGGnVn4fgY9umr/7cnsBLz9
NhO0VB0B1w5xXKUCWj27kWFT8P/L2VDPWF+p8BgjOfo6DZox+KKvVtrumnuMvfBnVq5janSVqzFh
mFYD3NXtCGyXiTRNkdHg9k8WyStGj2GDgGIiEdB5QHB5RWH+7PhhRnuHBiPJ/ZhngVrLflxpFM4e
C4F4gIZxvBwgNQigUv1m1AC54eouhyMiYQaFAeut2ST5/NSzKXjZHPpqY0sshsrRNkBCF5lNqWcT
WMWc0Ty01bytHTCu5HlzuUlCOmrNqT5mjhX4GC6OHgx5XhApW7PKu+csi2wkYKnO1Fq7fbM2HBdV
OBvAEVEJ46bHV/I=
`pragma protect end_protected

