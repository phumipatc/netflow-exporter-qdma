`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
QbKilqMlfBE0RgYIlZwfETzQAqbVyRvTX+FFgls8JNpKyi8pjJQwdNppq8mFtz2JhjfWps9Mwimb
bHNjEcmwx/G5jWkxIe9aYGhHNdsT3pyWVpQgVqilaKUES2ymRrhkUa3tY46tNr8tJSX74Vh21hzj
g8niJb1479srFQ1KBncLqH/TCYYM2Cf+Epjft4sk+1KtIieLHsl5XNBwfnLI9MTaeDQOJBHZQk7/
UM0D8zuR52ikI+D1FxWk2To/NaZQX3IBBabO1dk/d6NtM6nWl/ALWjvcqpK6bDG7v85rQFfYimbL
hEgYNyEDzu4oIiU2qcYZePTbPBob0LvLyle4EA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
BWvTN/MmRK+4hjPTfxrDD0gdItpNvWOom10IXcrGZcXNbo5FFKQGB70MSl8oB+FHNE+SXtcyzbXI
DWAMvPSt6TZvf3ZeXfEK+eLokJLFQDpWnPky3kuNTaA7mYp734ybm3sdz09sgQqyxhoIuvoa561i
m635WQqjx8Q94KLRoGot4NaeMlcRWw8GyznsxFRaddmwB3mUGXTVTkc7kxwsVqSYuo50siryDlk3
MB0qY8TQciFg5t0jL2N6VecxKsHT/MyVd9BmXOVdcx7j1nj/34Lzh82ra2rGWrRjjuUbvOJGKvrE
/3TCxftMOV96XqXi3IgYqdlVs99bgYcYSj9JpAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
PCQyEjN5oSdi/243Ffr+4dKnn1TlS3/IK3txtjVQmW/Jc6WUvfQ6MdDm/g2nHXtA74XGTEBQSLBr
kHL5TyuF7g==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
CM0SU73cOquR72ZTzzlmF5Z89TetpzYiKEX/+Jq2MYvv1/hTYNp1jR3LcIXmWksMP61UlrGgyTTs
4MyVSZQ77SuA009QgPdsn08ZB8wtZejxqyrg3X5agi1je/Jn0ZN2mJ6q2Rk8CTiIrOe6RsUbW0Gr
ua1gtY3FmwJICW8o0HFZxErrIAHOkTasqY+hKfOiwWqU5tJQ+lfSoWdkGBbNFCUVr7DMgqphz4u0
90mkzmaDu+YpkgvOJTPm5Mz74jmqGEo04AXbTKqh8YbjobumQg0n1eioLfQPmnNv3IUqTerRbxGW
6f0fmwPIW1yHsVNaJomz/nNg1xFJcAH5j4nqaQ==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ui2+/bga+1TSjBry+zvfZKNnDkyR9IPgMjgVXA5qZc0aDTU/S6bcWiuLzcp/c3dosOlG3RavAuUo
owyiNwYsA/R9Rjsj+pkojKCU+WLbT9Huym1UnSwqeJgXQ1Qtk7RIvkZJOBE9+1NQBU753aTvZFW1
ENvDuoz9gX4RkpiLywqbsu7VjjzIM8v+kKsCBsEIMtzny7bOcG2niFAEw7qA4/bnIVklYLU0NW+8
IqX/N6ZVyTtj14gzUT3OGGlWNlUr+dwwt8/jhJ8gncJu0HEQ8wB6KPACnbu1nsf1OVMf3OyHeVK1
RaxC02F5ifKnJKLfP9by1iWat+tL17VwlsorXA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
EQi74BbRXITdi2x2GnMWtGz41dbVufhOgdo2ygdV7qXq49P3w43buNQPGjTBqMYEmD5s89CSd9uA
NuSrhq3bqDNC9YEUdulmPvteN1SnGqTvD1Qi1j+K3JwNDuPzFhrGNhllhARhNLnk5UFRcOEoYQX5
Rh1TjCcmTT9EGMR1jE8=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
EajDsg0Y5RbzpDs9j3+ZFR3OBuVyo8CWsDLnYB8zMO/kfyafXm8Z74UUWHctTT3avKza9xa8e0dO
7EMwHuXh+DRdQVti9odUSPtcYhJp81JnfD4BU+P4/W5U6ftFQU1G6bPMOTrD28ENaJ0DzO7yZqQJ
xaz74+wLwV/ImfvndazDJZza8hnqjf/HU1gwSp0DGoVfrstZSUXGA4z9DWMFcjZ+tgoHPCRBcMtR
vBsjfI8zruUmjMheycvu5Ejn8pbq+r4qJtaooIy+8vZOhXSgylKoev5origknZxILp+upbL6fyM0
7ZTEwBCFwNHq6ma9GVTTlNc+9t0xqzRPccb6Zg==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kGlUZQ7DBDjUIQ7no4V2ZhTgfqSFzV6xMixUUq014TiSTf1R2HzB/KI2Z+RiOhVKB7+SQoxStbLO
Nbc68nxoZfPlol/HK4H94y0OcwKlXUMIKHXqOnt4s4qQZonhjROktiJgHDHP4C4wsTL61//owi+G
dQQY3VWI494+an5bKES9xOqLTB8cMvCO5LNgh/uoqrP6GRfcPbAV/Yi6IPvz9OiI7yv+5yf7z9aT
gqjF28K06f89j+PVt5NQOVEkzl5ME1zaEbT/ny1zMLsCC18iVE0XjZrYrgSkXFIgF/1su8ic89xN
LCP1OX9uRJCLAkW5l5Jwy0ySrkarIP6bCnp2yQ==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XJ4wVURF4JG9O4GXPxIuCXqeGa9I3i63FUp19q9XkU5gS+o4CPRJK5vUFqtTfaJoYOnuKyIKNSQK
YVcB3sIG+Yn385b00hlrGf6MHXWw6sCBrLAzAREbLLyoLyH54qM5/uMrdljnOLDABjMh0YeSxNfD
A9ma7JVL7bcM6L+0WGM=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J2DNDOegAKPzouW9ozOE2e0Y9dYettl0bstNzaoBOKQ0cxIz0ymlQtlaW8L2Hw/uZqaJ1P9Qk4Gu
uXTBhcHVB7mEBKDwu4nhckk1QOjCAL2McToitD3uU4qp67sjKYTDZBxkbFV1uaBwKk4IxvPVDml9
4CtKqnJpFqVDLvz2e65ufpzuizVNJzKDi+truSWXiMMSfi/HSqhQ7Nm7rO540buHzZaA/HneHCxD
HQ3t51q35mnDyZ3K3Ss6NHrDu4wzQGB6HBDXBGDYPkVTg32OVnv86AiY1qIJSPguFhS1kDG65xNc
vnE2jy7C+CfUjE9YW/XvC4S3Cysbwaqkp7vxtg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16816)
`pragma protect data_block
9NogEnDLbjyIs8FB72AJeypu+wEi31jdsTTVF3hgAqwJjlhBfNA5ymPMKRbpImsK/VcUDgjPesMC
8/A/sVyp7kRmNaq3SPpg+30DRRhbRhkIifaGxBDfYI2niiciQemhAfZHxXtNk2U/5J6vq6W456PT
gtJYM93zxb5wnXjeaMzc5Mab/dmcnV/Cz8yImr07GgOv246kZUlaRbY3DpVBFVMmMAyaLmLskN5P
g7fsiZd2hCapvi6UUBN3sRVlnW6YE7RKm1BIZsfR4lImw6FKWWNOXoT/QFl++2Ay+8VO9ttKs1JT
uYZcs+75u5Nk1NHKkWVY4txHn3Xq2YqPZEMlAj19QbzljQp6n0u4C5XajLWuw6AEWCROfBmN21C7
zoBXUkfi8ybAoDhfqCDPbF0y52AYnBVmIDUqNgIVySJEaBSL9PjFa9Yo9oknMKS5xon8um/+K4W5
FFBGWOIVGTUYaM1WA8hkgZwEmAO0gVdWNorlh6ftQA43mU20p1l6WA3fWHP3gsDEMgoUc3MJIIXd
uHoWTMS3nRJvYKlntoesy8GLjJ6//mm90aQ/TgEBhMUMFieH8B3L/U/N303m8FW9hBIBMzF1HYlJ
XZqBCH3Bv65tvTwpcqdeV+Zi4as9zqyaAc4Vf7d41B+ewsfDzEVuZL1AwahhMS8t2o2ruxwxGYSv
EMGb8TZZBzmDblvJZVILKXxWBdby1K+xczGIWkefqLV+2Av2TGtbCX4wDVa2m4gVWdEVBS9eeWCt
aU6f5DTbENUlxJCfmH7zo5uogch2d3NO9Wv8dxCq7TwYLXesjATFJidYYeTeHAjCZ/JmSLTECdF8
4QG41sRHiHmupkIhJsr0xFN2/6Fzdy+7iI9TOtSPMGN0bbGJcJp9vHw4BialgmWU41Jxo2w0httm
8cYaSiL4d11IE4bcbgwTqzzZz6hkDrah0gxYOd37DIS6YFucTWyz0OBThF8okl+BI+SUVz7t2Txb
zpHBW+FeSK2rIIUhmuv1RN85OGpdYJAulGC2PHpLzgr7FJ97vpUW/yile6uhfGv16LYvshx2UaW+
j7u7y9RTAoXyr+inkJGTsONcFujKCLtnH9rfECOTckw7k+7c1O1f+k/CBVpJfv+hJieF0ywuwcga
fSXBPX98hbXBPSvByU6PVxVzacCB+16JnwS/+KlqCStAUxt5S52nq5BadL+YCr//A3VSNdUGFNTc
dwqOL2ihdOW8CId1RapUseLazGlEq+2wFasToGorApVuzs6qh9rYIfUVAoRedLJ2Wzl9R7qV+dM8
5OfqEh5oN7bCS006M151cJldTAoDWJLcXppKIB44xb3gitdIiJfew2VEI8Pd2S1Dbl6dJ4HzgAd8
oyg/LTnX/dmQinBmeS48xgHMkEAVyYwWP/B9rya9H4Y7Oe+bZbwq2jqbagSFyk26vmgTwqJFSIWr
wkwh2mnclv6O1i81UW6KwHJOD1bj4cYthjPsqrn1afXI/3+L47PevAiYUv12A1DWtsXLzSVvvFdd
6nthIHKMb/E4Sbm//I3AywUxojI31CX5eKV3NO2JwtxPMHzFgERM4fwhdXMP99Kq9QIOhxrws2zW
SntFhuJkgSupqxwQDoqs6Pt3GY6/MoIpWDzVSbT58JPm8+d5R0Pt3+4OdVyxFVVQZRcpu7SyPxtZ
WuzPWtieOi8gBctb6R92PoMnLbJhu3MeJt3mtseoE0hnmy0YZ8GJeSXbXEJ53sjK8S7OlnyEaGkU
dyLrn+w3mrXi5pKRemcT/GBGo5K72b7glNFfix4l1AMujkliGNHrv+tWFM30GFOrcPJUyg/61dH+
l12uEI/fdK6jljh/hYIRuPVQU71cwrBGEk42XC9aJsQZ9ki6yMoi9eYFEmato984prlvDXRs/P+V
lHeUh3vdjHL9yi6+zKcE41SPOZ3W9nkpJfHmWk8ifwTg50FyZ7VF8ycig3YdxGchabZ/BagcCCwM
Y4dSO/wtiRX/4txYp6cRvL+VLw5vSElNUs9wEelQDm4cFqRzljmewWvgDIGN2KKeC9wQPZiy1u4V
E1n58lO1/IAsymQdXZK5zMNhrUysmXCDc5Zjt+j6ZeAm4UfB/LGCDzGLb1IdhuVKvXEjjO4KLfb3
Snk+rx3ytA1qir+9tzzEloDlzmFQ5YCzHNX74Y2ZNO06N2ja6mWPxTCfeDom3zdmJWoyzmazBghz
78/xrFk87utJCTucf4kETolskhWv1DxT+i1CUyqcw1al6qZ6vZGxV5EXihIeBCzysHxwxIc4IhAS
9qeFv2d0wOZonmNIPHu7RG+WOD9It10rG77XZQNBf54l/Pm9DnaVZGSguKqMJC2osP3E+UnmmJwB
27wbrgws3sdC+VWu67T99z1EWjRqzpm2bnYCvSfnK/mDq9NHkpY/rYJg4aFo9yk3Kil/qBkDOhZS
qNQTNgMu/E5e0QonBVh6FSZKj7m9AvOEP2iTIQF3FN7lc8BR9FWjSXgma94If677n7r93bqWkLIq
X3GswhREPrpVQYFtrTs/YtDL144dq+so+slHJnfK6nXjlpuXwpnPHUStBs/Bat5C1d61SDQzz5TD
mtM+dREsZIsSzavMPYkmvxfzcn4K5lSi5siR1IAB8NwzrHdcRWWk1EP+uTB3jhth0/bvQR8rCIIK
ilkY4iqQ66C7tze/0bIaWIzc/3Lo25bqXYHp6uEeWEzgfqS/Sm5tIQSKg6cx/j+SExYenprPVMm5
M6wWh4tVvjSTm3fDU09HznQNLvLBvEtQ2HUZLCSzb7JhGGrdmdMi4v5jIaEhCrr/wjLCvgXgmYZW
qBuFJGT+UiipdczlXcZTKhzgx3qil8vhxVhGkcatmG/hqD8HNSYc4hMG/6+9vFVQ3ZH4yNxMXdMh
WZ1agLBtYUSKdEf+MczvfW0TmhgKly10zu8oj9JyQGazpeT7MA6zMBbjC5cdaTAr2n7SVvYZnn79
n/DgDQnXzOrLYeZ6BbboHEfmVhZNc7eS1aNOYlhSucNlD1ozTJavvWEeIDnntWppIz9J22MkTuF7
oLo50tnE2DXlEpC57DDxs2owuPuaiHavPsyMJRVxbNLQK+9vVKDENE6Cd1FGtnqdN6W5QQ7Vd3hr
aKJEtfjsrK1cZ1pFvT46j+TbQPBdFjCKifTLIukNicEvkOlD3BsH476iGw1LsQhow7dLMSaaojZd
QRu0man5DF2Y5wYIHTMDT5DsI0x2FL1Gz166lkiEtFmTK9wHdxK8ISepgXpWQKcvCs/LOBOowDqB
cXRQgsWayTn/Hdlky2OSrj97AZFlUOl5awbnQAuNX5Ur7yOa1v39AIBwi5ku3XetGJ52Hz0Mmq1Q
SX9m1Bzx+HfYx5FtgegLja2i3wVHQM54+FWmTrQJyT4cg+aYx6/1tKl183o3btBYSE5IMNiKlME7
BvbG5k0GzxpcoiNZfNNSW5vFKJLJhG9HU3F+fv4jU9Jn60La11ZQNBiAabmOo7VIrSzeK47mLN6k
UT7F3r7vT6TP5pj62HDKa2UnPskc6wOWbB+fIMVOci9IZewfAJKIEI2P6xNdEyyoIXxfb6SqpDfp
8rokJWHXTUXJ0ZCLedY7hdB3q7/GYd1NnWa2hnL0uHpbY1bKEDeTsGCmbt5Y/KnqPMEsJFqX7MrV
Wv/wd2iIJQMA3Y55LAJWfPTCTSGZk/oExsjFcCVTCtxIv6LbZZtc4t8TQ9kp9NzAQ8/6annuZ/xX
pPbru6TIDiPPzUU3/vCIAXB55tZzw/Cd+P5so3JoPf556ek/Vu6LNv0GMJwbmLBNznjxGOkVtEpe
DQnUMEdOUsD7IGMFoSS02QOTWRjupuHysFfGvm25ospbq8YjbJkfoc5tjf/axDdxddB0g8af9CAo
G3B/gzfosfqJkDlkGiuirto5mB0kA2Z5WQR/tJJDvPa5hnFYn9xhDdtOHWDp3KHaKZ06NH86Ir/b
UnbgBYDiQVwSpo5mMYAV9vfdZqeKGSB6y3wCwCZrl/pdgb+Db3lzzH8GuRJSJ4UZsXk4Pml8GgVO
JNDaFkj3y1YeFmrbuz6gS/3gMumpqXsR72Z+uXTXU0kjf3qyujx3GN0KM5FFuexh3uYrf0ffVJvQ
445HJJHuKmO51BeG935btYM8odeazrnMFT9jZILpnwv73HdJd1cf9tstTIZpp6btfDYc5G8zE82R
pHxAmdlCG1GqbVpX0KuVf2zS2f+fsX6env9Q2xSRUunzVxadHrtIQRg8wdAi/Qfa58O4qthOcg4s
9y0433BwPmiALoYJfln2T4EDhVa4+hPrkH9Amu8ahQEPDUe2ohoFSElMGSlZrR7oabvgXeRLKK82
J6e63zpkd/jZKYF/xaMDmpiLwc5rFtEQ+cvrkl5hozz1S1WlYXmhADk+29OPqruLoJ87QbTE3VEB
4M7JeH4oOyBwIOyGfFnJRZ6PJXgKpnSFVeasw4y6h7JnU78naquwiCapywLBjyMDUnk1zuVpieD8
SMFY0zNKffoQ7TcPDf7YlwOWbngyFkd/h+tfQsBVVikmFd6Z5QqPhBUhkCrieCluBK1UIWac3d1g
k21AGO5soFTfBQxpHB7ekVbjSBeEyBmKMsbT92CJ44iejm+6PPNiFibANyWCmXfZOGYQv+YgUy9G
41zBZ0L3Im16/FmQkbZCXKb9gieo/sIW44wkt/fZjW7reSm/mtqvoiDb2ba7u+UrpPGm+hfdyYsf
rN83sIHZRLdN9bUBh6KUztOyq4mrECgnCSVUulFdLrs29wm5/SjF9eA/wKE0mhPBxqpxcRFa8rwe
eg458pFohzbq+0SGAqt3V3Co+12fzkMtJRmwqd409Fxk1KZGXFW63vzfznQd8sEUbm3o8vv96r0K
IAHBgvxB6MPHSMDrdJ+B7zyTyLCUR+98luXwQrldffjDOCExGuqWoKclTWbiZPTyjoeAZTXeU1tf
A+NeZZQj38jxuyEB0O2mt12jaUDQk4hdkfdhGVbIAgfc1tFQjfhh8ECDPW37LPvo0XBQTNMeMmpp
5xHsBdCCPf2hwh+t8AsY4E8WMqvkce1ijmqMk/q1NKmbYZ1En/M9341f0M41vZlS6c5/1YJ3h3Ov
4PJq4RpCOkFiEu74E334ZJjp0ZpKlH9kO15GiyWyxWIsgtCMmTRFN+FwVV+3QpxiMnB062EEyDrc
9e1sGSGIpNdj2IFz9zNhupPI7zX3AkMc35ys8scJ7VA9mcJ/ebv4Px8Stb29G0ky1tWDRQprE8Y8
akrLfirgk0nQuNLrLl/Ho/f3Fkdsq0zDkAcLVTxwZ0Jywi5IeJAAOcre02z8rWIaQIcDULmyipIZ
9sJ7QY0l82G+qFWSOCN8ffr1G/CsiJJyCdhTO21OzrE9oPh9PMycMHAkRaDGKZUYmVPFBK9LruLL
PKlEptbPwvm2TxcZvQwyNOKw5MespFXHO4NQTNgeCQq4TaZxf/cFW46VrgVJVQjrZntcr/SWXeAK
UXwnJlk9QRbqXmRz7CwZfYTCM3mMYPdphpca3vnZ2v/RvDtTIhZIruiQ4BSmbyOVVNoNm1alc60U
0HTZMyamJbx7YSC/rbdFuhMmB5KbMmuljC3ckAs1UBLPFeqFyhQ/BSV1NTgcuH9BWmhcUUR+sVe3
0/0Zyen+PmOPjZr2cTzP+kkVhjd58CbpSh7rMNc/1piVHld/qIukv55rTX8K60xCr7wW4ccG+fBM
CpsNQXXP4yE6IRE8CE2rUI1gXgqTbb6ZVXpYt9KfS289YFr93xjBJapLqmMlY8LWlRGKwpx7v5hk
Rx6jip53p4MgT5v3nnj2YJSgsm16LU4AwHW1B6G9imBEz5wZxoGo6xdev3Ch6ydD+zczOjjzyzB0
AETUEUiEJH8MngbN0R1G8B9JGE4DoVsMxWn+y9M1/3CpMHpodnJt4JuzrjOqfcIPNS27OdYBL387
0bJ5hEemQZgjX/7D3qWhpuQAr86O4JPJkqBA/SwafrYWt3KKfjvgKF2381zRjiNp8Wwmm6WNpO5W
I/bM/Yqz2mrtbYVk3+a9fnAuNQVEtqoLltGuTUNWlQP5pIzFOIaaEqH0C9+f8SMD7/0BE4WXrbvv
ax+BYjMxTkgYM5PoZ7lKqZl4BUPRWy2ZnGlL8H3eCAJRAE1F1pEgqdwPXOkHHGu94ULoMH+ZfbKM
l2/S70R5rd3cdKI8s7L/yKghJ7KyHLMCVJDAtmJuE3kJaG5C8AYXStPBlrXLXlCZKLxd3dsRqD4q
n8RlzWBHDEa14F/Ep+oSzfnHFpu2s+KudA0MIygcrfk22EVr4VJpd3fQZcY0Ca74hLyMe/2Ec0Uy
z0sHutrmRei7quynT6iKkUHzuP44AOa6af+xcVkrfEtA9Efz/ISx+83PdQjgOIPRMr2ZvW43NVyj
6Viyl/Nrf5uIIiww9j/xA4iPOPuZzO75Nz1TM5xLlMzZ30Gk+5voJiJVNLCJJYmduL/dHLbwx9bi
2udzIC5ewzlBu682yrGT4b4LHVrqweWOB8NVFlid69I/enJkg36loH4dYpuVRQ4AspMeRggcT39c
hlpkXPxJLhvDWDnJ9g9rxcccuBnL0KXT0jA8WPO9NZL2izbil2W0EdHfWue5D790ytEvJpWOI8cy
G3RwTs1PmReHkZk+Aonp+CZFKHL5hz2GbdD8W8/o43iiW39JtSKImzUitmzDKavBeN2CUT0cNUy0
Ce1fP9b08V8qzKQ+C7SRfwSE3dB5r/li6ZgpYGPbDZsAIVbah6c1P1dtN1p05WWKuFvHCpaok7r/
ekEak0hIIUoCRbBDEmJa7Dl/5M8IbTbLY0UUfkT0pegkXz9pCteuA9QOXMTMNhYAuIFjEfUO8Rai
p+FqlqrjGbtHfIHx0zKpoaF4Qg+Kgc2WeYBFqx4rC/YG6nuIiH13QpNz3LAu/bGDRKpW6ojHN2er
AS0mhJRWC26Zo0GoY8vv7gsR4TfcXtUhkDrjo60sLu83xgtqFT/68AKLz6BKAbsGw6guMhJ9CLSK
5ify/Xa1V8J+Q3QW4cvucXWjuBjH+6p0qHFKWa0hdmNLY86m9+1SHhDK3gdzRyt4TCx5XiWcdZXb
kzqrbqsNzlbge+b7hz8XHLogDtlydbrFRuUQK2zIsO7q5F2D8vierezwC4DY0DxOXUzC7/Cgkcvc
NB+v0INhsQORmPajGFK7E2psiY5IPakRHQfTf9pL73dSLZP+EUpYyZAZP+7sd2oQg4uaeN+IrQOg
kQ8d41jz9s4Y8qaYUIPpOsl+R2Ab85EELRqvXQjlmBvIDNrVuWv626tpExR8KAIlcDPA0ikA5Euk
Wuoj8JWQQtn9ERlOZDPxJZmU1epLoeshY7iRqb67HHxBkKyJzWYDGeCjq+KZAd8EnpR4dOX6lddp
0mu4qAgyCzVtjjKRGOoui36/RyzwkYaNR6sK00W7FqLtqoBwbym4fHSNSKD1DHMFlWfNrz6rbE0o
OI8cEQaslan2uYpMWAFdtKLAbsnfH2SJnIhLiMIv0MMkPB51DVGJJlcuPZyBz2/iTq+P/r7I4/nz
F3+xHy/gMlw/zAKRWLN3fhKOho1hxWLDq6dfdHWHdqtViEUub0kF/UGHg84BMCQrM7jtYlmFOMTr
6SwVjKVrz182mwb3kTpJzuVsydR8xxa5VkitnNRXD2duaQtQkUXlqF9uYQsqqvjIg6pJdffmaRXE
NpbCRzy4Btw3yCeJyTAdW4TsICepvPEsEWOSzXA+GKW5iEApeylHGEg1tQNaBY9DmzVrpcC3EILY
b6AgM8Hqu5veU5Ls+SCkQkmCEncaDRkCfcavVSxDqmVK7KK434Q7WcD9EADkGTi0YEP3fqL494Wj
EuzmVZdFTyOH6OojdFSlZSKo4XDf44G1jr32fm7asZASnxBwFTVObtNqCZVvOhub1QYrienAIjtC
FkmdtvWD6Aut90ppaFm+nbH3XcVBKJ9wDzq33mKg4RDvJunkCvuFxhtA29/We5c3YmR5MWzjzmQz
wUS+dq3tKbp3/RJzlol8nVV7ZIN4Lzp4B5uk9V8e0f8G4/lKcMk3LbfALxzNuoDijshY2++f9p3U
DgLmqijjOZrKyxoG9JFbGsxXdDIOWpx0Lqg0LsrhG/zatALAx5Vup9BtDdUjvFwq2Bc8Z9FmR2KD
VM74uReMwLrwrebhPzQUAyz1tw+qYdyiwgX7leqvMFUWXELqAkOEjD++ixiqdT/NgDL+Rm5sn9it
rYiDO2WZlbmNRTPS1kYBl5FY5H6Rlm7T4nMPH9o2JmUEwk5gCZuReeqvIMlBYI2B06XYuQZRQiTi
Q4kHbq+0FLyO+PGRtk7EclXBMX+M9bHdizURBZOn6p+qFIBZFxl+Nrvtx+KYx4DS8qdSmT0m0Gkf
OimwJgfS90i9iWfiD20AsGgyNd+Fb/EqNksrMhbmoiAYEwO7bFwBVq2p5NxasyC3/K35HwCNaraQ
CUYQEMJaq/j2459mrPXii/lvrup1LOk8+SJ2CRoGbi0bFirFF7yjzJwBKm8A6rYdI2cH61n1xDTA
D5+Pqqy/yX3sezM3UI4JvdIv9WdeRDF6keFt7VEoFN5UFZAPPRyx8KAOYkzMK9E/ndyj/3Rg+HFj
RGgSPaBxc7JBPf0fvsYpUKPMJPHu03bC1SdGLdJlYCWhqSAnOF6XfmeKWlK7BBB9/aBi/AYL/V3/
V0BloDjVdTMDYcdA/trf3WhHdLgYifLiwOCXa9KDzwz9irvpKJW3gWU21S1ABhi9XvW1yoGOAmpz
2+xVLDGId0WJ3iZgcGlD0lsmtCgCfoF30WfrSVh9+6UUiWAG0HLwH0j6f3O3t1HbJ3YWAh9766s/
MAALXmXGqIkyH+EavAlNv51IyT6lEYsLH38p5A1xXR61TV/3TLmYGKZczjyGKpTQ8V5TfOP10bFE
qcevqjH2iYes5GX1KJXH8SHNSm7lx9PzuMr/jSyd/SDWgySTeIEAuXhEr1Mcob3Dati7jyXxKkse
uuWm9u4+vSY0LYarGB2f/ZnwaIe/TRgdOpRd3WA2UjxgR+sUnVGVtkUVfzqkM1RFnQQyFMRbiY7v
rwDR+BKc8ih4ZRq0LSI3UnRR9Wu+6y2fbyp+T7JDONPFrhepIiPo0cmoEEQiPaIrteA0av4RIYW3
gDM8mxmMUaJ48gn/adDH6I5kjbX/yaigI+eGuSo5N70dpfBuI3tegKy+CZTWFmhkp+HYBDwOIbyW
ycPoK7g/aRFboMb4p+tyhAtq9x+0AydBWx8ESKIr17kARJm/9nMBEG5iXMEcMlYly+8jXMMPrI2H
jCfMLX/pDZnagk0Fg49n529lQMAA/Zd/CmnDFRvPQTEsztrhExg7rAy3L6V8TuuSHGjMUUnEXjQ4
cQszdnVZa2Reh+J7lvvibi8gOutqPMaHs46Cs7ubb1SGi82RLufyivrZmoYLUBAy7v6S6pKJdn+i
Sdptj+nAmsFT86CoQ9x4Z4cnMnxEM+emmbnMGK9xBEygQQ/xbo+lgmo4buvQD+hJE7I/tM8kQjiB
Oa0Rjug6aybU4xIZgTNfBFNQ61aa74lK80kIyNvL4cY2uneQai8lFiKAZ9ZB4qIViw43BalUqTE+
LIgmrP8R8PlEDPxWJJdM3nIAGfbQdW9jXQq/IhE3Ufvh7sJzAdoMW45EBz2/itI9F4LPTgVOcQRx
SG7nx2EYcp8PuoxZYTp4Alia3f508VVNScUlvmRrg/01Wl+Gi2devdqzyEAhs2pbt3X/49azWtqP
082rInaHo3KxUruq9Ixiwdt0QXq3A0DseBfLRoyTHUzTGY7Ba9kRo/wKsRYApfJIHEXMRMOc0qgs
Vhsdg2EjuK/Mrp6XNBgGods49KJPZ15fvpxwmFjxK8vaxXsoyOs6pl4ctZloAe54x8UPbUvNGG4u
zlYi14p+SeG39I0gCDlUiOU39hi+rgFTaRPXUuHTKwA8E0b5NIWhG4AeXs5NlX4oyXXnPW4vK7FJ
Ug93k6XaGRIKi/GTrSFBy7TZnUt+1NLCSf32PTNCjYP+2V51WOqOqfmIiBkhicozPdHhL75Vw7Qa
BqU6/jNL9dro05jbGCejuDcIjS8Kdi7K4ShyhsmiqzIQwDYzTOu1WkskBQVC2TnT0JtPL91gsxU/
2I+yMwK226Q7YlXOAvizvz2BFRGl8VCDA5jCbomU1ZKv1zJxA/JSwZXHjKbzZE4PL3jqnH69tLVT
JhnvrPleJqRPPSI9jIp1R5nyuYctD93H24rr/ftGXTSJiM93/B2nQXAVafrj0svMQ4SmLyP9yyG1
/CTfF7VNH96GLNGLxjQhjFlbehaOY2Lkr4yzufTQaUV46rJH9sOS1f+hSEv4CXQDAfiFETfPVjCy
XzW33mbaOTF1c7hWUCr/aBwEu39WeZjsRutIeQy97w4d+3TirQwFmBVoOqt1J8CBH/3RTCA3s9mn
hRbhoUSnD59uqYh7PRYYajFz6CNW0krExGavRiNw+U6n3YFv3IV/FgGhLrohE84FvTMCbW9re0Rc
7KAhzxz34KXkfdGKmMBpaTuyyvWVTI9eMuqjVVs4o9SBWs3FkGm4y4Rp5nzQ1w+xJkayxnJ7eRBV
9GglQMoF5y+uI5tEZ99bJ88bEOJV7iGLVDKNeuE4Co3Qw8NahNF1XUKFnAnI8fuoOLmB34lpdkpI
wIWRULtHtzZDlhwRVLa2GFS5q0y31LGPmlha+RTCnjQ+GzTbQkNRA/EJyVVcrYy/kWWgpQ+KhaVT
7T+vATWGEn6aDiV2P9PF+SvvTsbXESUesyNpBiTec+LaYoY6tfN9f2tUa//8YOosHZPZ+/tivb/T
ZZRT9ASv+J/S1UNtD6FeAOES3Mf/ulhq0xhZnRc9fZo6i6z0M95vetyJFZ49F5gbVvJfqp6pbIZK
oQ2aykvnRo1HRdYQrnHVXyT0KF/ImSfkZr6vWt+iJ0wFUzG+wVaiwSgIpTMRVgAO8HTbfXZYsTdM
DcKYfGLQBaF9dWMJu8nQMl9z1bpYyQ/iZZmMx0V7lt0Zztm20zuqMKKYUGNuK3qe7XBp5E/Obf2L
sOjnFx6SdWRMXtPsV1Cmwht8l2CunfTuFy5Bf3K9FiMur6X1RIkXZVEB1sibOgnUvusdlKJUq5Ip
/e8Tfij+MSvzcZ/ly4I+e5gmD1uRf3uf8syfIo/OCDRu+WEvBiFJCJ0pMCjh5BfJlAHroWGag/H4
eSRd5GE11Q9uWiSQCobZI/YRMDNFlaSImdGZHgodWhaXOFPv1AC/jozF5cGNZn38TmX24vrY/8yF
PjTb1+tPM8lgXs29cebXdErx38pZ133GPiGREKd+lFjYMh3aHOcD+Hl1mvaUcKkCuKmwA+zv8j5d
hxPcP65AXPIN3CtVzuV8EQmQUQlaFVAXWG+SeQC9kxhik7ds3mMAXOEEfUOwpJK8dUiferADMqSW
2yXksoGRr9oNtNUwHyAkacpa4/EKeFLf/W1vDYVqt/tePaq1qf+vYokGKXdpEi4QJKKNcHi7jAVS
nJGNjRni39EUakNfR7RSPmf15VfLct4Htl2KgDMhUHvUuJNm5wsgM1WsZwqf6daD0seOdIW0oYOJ
7jp+XLjHiY6I38A7AjUcYi1hoag9pqTHkC/noQW4iVvUJ9AZW0zbpKWXUBbISCX0fmfb1z6zkTvJ
zMQDVEK2OdJ1iDpwDMeqViYRVLlVhIiHYq3hclw/EilKDbJILUWDKFhHUlvfzPfZmhjCKo7ri5s5
qxzdaDwuuzzeVlyC14YkfUmeCAoSAIxIsOHc1D/zDXtEdZWVQn5unTUmC9qFSrpsSjPOFQhs2dYy
old+yHWfQmL4ezoHQx7q9ThE1jZibTTAut+23sRu5tPvsYWPfN8z0e8elL75ZmMg/jT7MLJiRiN9
P3i4r3SLF1RYSmXf0ASQOCgcykGw9250DviL4q0hT3399tX3png9ppk58HbNnXchvss52Tg/Jwma
VfY7z2zD5EHOfr16CQciEz4PPyLGFd80hkuJ+PBLO5nNg227zwPAxp6JV7RMZt1tSfim5l+IqgSs
s4iTSvzmlSy8HKM2Z2naj+Bny8PF182BS/I+sTLMYkn/M1/F9Iys0q/9ZnwxhE7vdJZM+VoU0EwT
Jlus06hr/8Y64AtzoReFK2htm4mKpRE0Yra0m/4xecmu6ckxSF9eLidxoY46mteJfr8vvSujdEk+
tdnu59WsKi4wES3BIdCNkM4NZwTpbK1sJYaY80J15WsNNtlvfXsz6W8UrqommvpObNJOOsGkb1DR
lpwCcLPOKBTiZxAztbawIWathTSGBZsqcHtsq5igJ/OwziMPkmCwuOOh/8ABtOAoChQmxPg+J7p8
5TeLsrpdZHC/3aqXo2ySRRnJUEtfi6E5diLVMJR5NI6uT2bCh19WaDuhM91nYr5llP+9gd4yuUa8
vj936o1tD20eOGkGV3vLBvq+UFv+zl88ktWNiMVS7vWge9SKPrGGgMUrp65NN1yJTRIlQnnMNJal
4LoqlSrVmABgd7NgnIRGyv4InRkR9Y3jl/2xJ1xv7rocv/9iDUnmduRrum1xM6ypfezMRecAQoU/
Cj0zE6p3wuC7XHcfKTmh0WF+kLEZ+8IiYzBkMbVww0Nk26zw2/MIewI3demxx8wcjmsLm9P5sswD
HwDsYSik6HOfh3qOp7pmEtvZuv9t3P6vtM8WsPPC3rNAld4te01qmSkOfD8IikHI3NwAI2rsQYt+
sMePaC3Sp1o0XTjpUPsPUjr8IpVoQfZgZWni7h2c2+rJCWxOqmN8CsR++FmbDfFy7qvDaNyVk4aX
OacxjB8APGMz3abJdSdZaWLbanvEI8fCkGnmBpxJOnqBe3PtrKb9t352ZOskhhC3OLnB9lh+wrnH
gJup8iFHWCsBtb+o3rQEQ2lKIG/XYd1l30IjhZVPG+lVOBCL4WmqfKkYWFnXRcni0NPuyeyINNHk
WPZLLAnsdWqv5OZAiMzmJK7amj410up+emLrdA7Qu+Y8goHxfAQqs9Z8Vh4psWjtQ9Ht2xKUTo7n
YDyoJDx0qj0zepfVVd2c2ijV87fT+dZUzYqsUyliN/yUAOLdbmKw/dgJuVIvXSamVqQA1v1PCncJ
xUcnBREZjSV9dwQb/4XMe9RYiWtU+fG9MFpEzHgxvGQ7vc/3bgeiWKdlQQNwnNTCRCQ8soHxEzA4
7YRH65lqt9XhfxLVklm5bKyrgm3mqAySpFhiRw5jzr/1aVE6kP4xM4q9hb5fJmgCp6MyIJ8lEzON
pEi4duonVPWcvSTaZIqyvT1ioLAFagHS7s2MhNEsIXVes+OQ6cYAthSCPpGyAnGxam65Dh9B5gQo
0ccFIH7Yo/kZx0+wuLBxLcotzEeCkD4WRc0G3I+d6UAtscto4M6Wxy02L/wgJDnreyWsxx1YG0Vv
2r8G4fBTApDLm471Bd/sg/VhHYDezcKVoUECXSzt7HCWqdgulJGiadgcSqevoBj7JGEhL3wSi64+
q/zsGf5J7GHMCwLiTnBz7i8pyu7pV1qcZwOZpZy8aF7X4jaT5c5odf9B88kq8KKtnZNSxWcZRFGR
3J/FaoBntoP/mistIGgeqxRw+mchbPfuXVsduyUegEd+n2a5uKuoK11KVtHRq8WtyFCLQSUrZPdX
qjiMnM22XlDePGSW33tm+AB/E7cPOT8R7mTMKqUzDaGk41LYxzWBdz1YaOSGxELRjTWSwRbC7B8z
LfSUaZnIynRKbCcSLwXIp3d54iXQ2k3JSS+Z1Jk10U8BMxU4L8E2g+J+cyV5rVFFpyexs16yONkM
OSeaXbQmI2ATKv7tyHnsiwxOy+E3ZO91e3KieNxj6aDiJUYruDyn+6y1oHo4D9pMXP+cz0HfR1lE
Em12WwXJhR8fpv34IDsdvsR96bvKYIVC5WBYtcY802mtMiYTcL8oQ2VpA+idgEiWwXQGbPaP9MuW
z+z15q3VcoNRl6ECP9OHOtwcOZ8GjzBgMfe0hdfCpiS/4/m/RvQ7hY7ZfVhZVJ5o7ZL8DF3aFOHT
jzKipmrvzYu/WKeeDhomHV7YWmTMbn/MEVGyRT7xsSqqwOIf56Hh04jhghrN45dJGwaw1RAh//UQ
2HpEpVZzOH6/IEuUKgkM12ItZOYH6qlIoFy+JlrYxcQWkq8YS27BakImD0kDm013VqWP4hDaUZ0x
4mbdEw4fbYemdJMfFIbS8mopf2uF8GpVXTz1rM3CAX+hFW4JW6PeDg/MKXF+gIzsYcAA7Dzd9whu
5f5rpOAWQ5+EGcTrr9+Go0h+StYC2adFtOaRJJLFlVPMPvfq80XUtJp/tNBQxR1bS6yzs7q7hEWy
y+7nC89BGdjkcSJeYzUWqZ5hxKju8/cogMHG/sck73/36+rmsdH6PG3YY9oTKDhHngcL1J06aL6/
b7OwH+uFqwf9NKb4PqG0LTrhKK1vsjnHMZIJo0+Lc0M9pcXNkSLrbgfs3OUu8EGbAO3xk9IKNp4N
Uo6z6DbH7EmkntKPIygu1i8LJF/eRpy/6a+5ESNpxbRXG325dww3FufTAGFxnprDyqLXEnwkRuqp
d5r+gmYfKnWKMB6jxClwdGg+AjmMECTgz8+3PCZMlBcVZLZt+mgZA+A3/IJ/cxQmhnSXeTSuEPbL
2mFPan5zmT4U5VD9lsXoiJq4KewJdUwZyUgLPk/ILPc5VivP2ZutiSjmeHf5UK7Du8vy/A2QyORf
XfA/QKEFKIjcxtBOgpunVjpn1VKqCYPY1nxex1J0l7XD9/aVsNyX6y5q3q/kuuIMVj1W8i6pVFdH
c3mZ6mVLOvyaManNOFa43jLGlsf8GcjAcbs7XoyubZMTVsJ7ckuo6Oa7MGPBCoZukI0ewyajfvhP
vUSyVnvz6EDCyGw75OBKnJ2wAutymI/x2EGUgwJAlvsM+1+hV7E8Nw0hfdjmgWm3gpLGbv7dXPvj
3HuIyqI+iRe4n+K3WsOgstZNaGiyHulTi6pN4B9lnG7qGj5XoOB7RH5tdfpoI9evE1jhOtPBftMn
o4xjMRS7jxUP3d/ZIrNmOV2Ebv2xNPFabGBVJAWK3OhcFEjEub/qD+OIc3eumV7fltzMOJ4kPdtc
pXds8KmBfa+dPUIhvw3JCjQpHMeKafqPJlJcQjevmNBqQba3c2bTrHF7VP97zVRDv8+Z0FS9I2l4
P+214jKytCiaW+H4qpB7VRp4gmuiIPEzRTswd1Iw0hL0Pk+9g5Qhy5sl/j9QZHeTCMj7OtFlCOMe
qmGLjn2X2uwGvqiolifIYJ+pLed7hfU/WkaY1oaxeHFXEIuCKWNBX3Tmfiw0qZzuwaKl+XaFjlJF
+V+//iicLfos54PpITnU8C2Ha/1ZGkyUJdAdP4Eb1Aar9FI2soI6JqWf8W16MwlCtmOSsK3GpCKO
OCYPQymvxjlVP5H1ql1p/d2KlSGY5on9PynSpuOM5I4p8Go24bjELnu0Ip3AQwq9Apsaz1r7C4Xn
WnUP2DfUFQdX6Hlb/jMi3tB5i8imoG7r9/YSOkuiQhz9AKD0aalXiaoT4p2ROr7vGZioltJOqKIN
GxnFkLyD1zJFBMvCouQQ5sY5b286d3aNwwRq4hdLQo+9zqgok3SYBK9m4pvqF4IRGxln0p6O5+xv
HKydPpyA8hswBLc5FSVopToZEPDyu/ekX5+yzf6E3+bacF6ks5ooU+PkXaqocvNq+oeXZUr7W8Ve
3CgxGKQUyutgcs9jXZiPZyZCjJ/cgDMaq0tbHc5ofmnyrLq4M/RqADSfoUuTGnrMZIFhXBfH2syX
w2zPfnshxrt1MAFQpUJ9qORCOrxhGr8ao/h3SECBwnc5Huc9Is/TbydVsTSzd1PaSvKutjmONpX4
/HKYi1e5HR/TPv3bFMY3ucRRByYbmte12af4Vh5zdG1bdlONaWhbMBV9Mk4iD0asA30n4S+j3FsV
bzmtHlkXoa+IZcuzpH1cH29Yh8+QiQ+QkUrzjaM7lww+GFqNJQQBWg9uXOWhT3MONqQpmpQZtu4I
9V8BiWxziB7jEV3Z/BelA1tWxKTYsjWgpJT12pLGN7ZG1AUolHOIzyI1c5Tf0Epl5NIrIOsAv6qF
Ex3Jqo6f/weWPd60Kaigjl+kh8mMVH6fyqssj6wrK6EyRQ5ZoPUjGzgdyBgg3h9JP1RSNajpXbBc
U6AhMdmtCrhfEEBiQ1n80KVsXua/TfeSnK/j34fFxZC9+Nhw63Hd2HK+BGYzg0eY8b2qGFhZynMR
819IQsr1xX8NUfnOuO0GT1Dih4dvFt0Ti4/CvBEHUvzlBt5SpfLsYA7NWRCMv86td1O5DTLkfIOs
bq1Gm6luil3QZueX6SU5f2eNV+GG+JiimIVBSj5UTY6IrKlkil+o359T4ahdwpo3Q9X2B9+MZF7z
Wy41vGjkpqEnAZa7zqbi/pzuKed20OnnIbr7hYW7bw3rmwm3Kao80ZaG3xrRNDh3dF2gchXsppKL
CR1PEi52MmWnKxiLAiHOb448szWkeIHEl3jGJwWlPaiqo+LsSRzVP+vxypnetuKocyvlclBDi6V3
E8P8Tkz9s//uIuUkPe/woHRVzwdlKGtJ+O2veFtlYVenmUehP9h5MvJo60al9X/yQ7H/cY7sNWI2
olJyoJaGxBBm2dWFc1gT01MGbbO8WNnN3zYAXc8xFyjy5MWD1WMCa2+mpxOnfAt1Y+sBCMuHf3c9
5v564Pm5GwUaKVskNI2+w9ZKz6jJ54RN0q2c97a8ZFmijxsYHp2g1qH/Mv0U1bS6GT+SvKPXoXDF
MHRcwOAtKfcbM8IfqVZSyRpt5/4iAYJeZEmAJnyl9QbeYhqJEgQAkEVYoRkbfnlNXyzzMNjJh7q3
kBCPMqY5E+3RzJofjqKbtQ2Rp+w9dVHwnWxdcVMFpYzFvW1DLdgQfAkQ/ynDC1RvCoIXv9IseioS
Qw/d9sVT/A7BKw+C2UGlDonS+Jy7rdpthxsAD467jlcoE4qsChtEtTmg3x1Nk6AFmgI1sgZdH6jm
9L1fS1d8g3dLcfe54y65XpplCoemdxa82f3fkHhljaD1L4s6dMrIbUoFqis8GkdWkENwtLK02+Cy
TUyB/VVlZEdelswllsCFM5yjTxq2zV4UR7pu6vBo2pdr4hUcC9CxtsdtJ5ETr/qpsFez1WVYvKFT
d8SnbxIjuEJFNg7kCxBwmglYBB3pz2jAlASt8ACN1cKK/Qaahl2BLuv5Li28SFwFsCFywx+jkRo2
vR3FN0FTmJuNeShWvEwSCFxNtDztF6DersAVJCg6Q8OdecqHeZEtp8NelYWXNyrVWGMm6VJbbU9I
AQ3HBJI7Ea4ybG/3cqshgj7Nkp/lJjFVye523uvc3TtnU3TqPHo29xnL32x9cOtjGOnuEL59BLyc
dlqnrv5gRi8CdhaZ2TfiMXqhVEYyNFXIBkykdC6G7x2HDA+ve5s40QEna3DzAxrGC+U5x/qFxdpW
aTPZ2qihWJeMqArpfxFuFrQDoUks4fhMvg8FZD18c3509tFiY8/2EqB4aoG1d1G21mqB6l+dugih
0A3oX6gXLGug1GLyF8WKapIyzkgkJSxj1A/3z2JdPxrypDK1bnFNW+yxFvPn/i8MH//JSC13fFIN
9IBog/3oYpXPZfcQbtpIKioM0xUF06ZO3xcgglqqG2AbCqfcU0/yek/Ik7r2lrJsaSN0cPSi9IbB
ZrsM8KNwlyYxTYRoQHIWdHmcuVdnAjI9OD0IXyJgJizUqU4fb9wUKqVdYRhxCDyMXczKQ7BvNeww
r90tR1LEW8uX4psjLmAQxWtk0WkyEJE7IDSeHALdDPdDgYzLoZYRvoXxn0LtheD0K4tpdXJvUOwo
hMPB8d4cHIHDrw98aGiQ/3PpqugzQ+7pq2cjrkc4ejRP2oO28SG3txU+4Qyv1SgDGHY9Q13NBMvK
znC5pXpZo3cy42Ln92iHTwXrS8Eos52lLrBEkjKX91JSztqynnu8fidJFUXNDDPW333HlV3j+od+
0dI+dHt0/5y85htzfcFOKtNjBNP2WXNcUdfXO23H2UmEU9m+EjVrEE7Mk87ixynaxOh5dxXLMc0G
WUfJC5P5nfufX/9ZZcTelOxqeUyUSQzRru969D9Ij5csG8M3uBMYOb5tnyAJU0vdFn6SyEG7ciBs
7UM0Vjzb+dE1dd1BMB7UNIofrBbfBzFQG/+4lDnneHkfWXsFPuWDnbsd3Tgpbx+ZThUyWVw5TAf9
6LgJ9mADIF2DDXSL+SbSSyPDjWv8FMf61AlRSk8Szi+gJMEDsvrZbJNMXqYhu3na/hra/iZ6W1U9
TGiTKlt2gJ0xVc1mqWuvXF9uQWIF4o21UEiYc0hNjb6/MfGMl19BQgKorhVcShSctPeClBynXh00
rF9w+ue0FchTxmTA/RyZPsB0MZT4lz84OIvpjWn/2b/4kuMFYgUuU0cZYZO0lr2NtDv3QzmaR3yo
7PzWU0M+MsFPUlkHu9CS5XBw8iJuYBYtp1sJkR6mKctG1yQVdIz6kIoO9qekQvYZissogPhzfwV4
P5ntZtYQ2F+ZUof1vka0NcO5vO2OceTip0/PL/t6gA6Y0DpF9wXrk1C71esXLTEotk620sbVa9w3
33xO6xkzd0O5W0WE4DChZVn4uh0euKi3hWazct0R0onsOFwJoK1ycrYH7FLFVIm+GoUdRMSKI7MD
m4UIif5aFTAZn19oK8W4hORhpHgvMjXRHhMnIFMI6+IT0EpZlynUShninUcMamHsgYvW8YbuuBjv
1NlO7vcAWbGtZXwRx230tcoK8ZpI3MkJ3uCjM7ZFgbV5HJy7iOUpbVav9hA+uSsxScIGYBGbdlSz
EzNNpwhwquCnZ0zDMs0J+mP/F7Yz2xwbv1di+EhqqSAaeZQDZhhwWLXw+uWI3sWcUj4xpBNxb8BI
ry5Gmnp9Buc+oJhKRagQyCZ7FqILav6D+WFMjnw2YgOUBo/JfOtVepoVWmDKmLCpaEupStazFTw2
Cz52b3KYzDocC1rw/wtSvzKzh2vO214vXIf3hn5BeVe/sEz9hlBm67rYXLUspOCY8L9rPxgpMsI7
UBZ0Ni9y5NEaCbbAtC+6kYd/VOMoPIHAKmYAqnmjrXzpQVymwX9QnWI5QNq9R4YQMWiqFTdoCSRj
FszFtm014je7BGIYdzVI57wE3mM4P3E61HS0BKq7Q1rF9VF+1FNJRv8NaGFbyk9KxIacg3u2bCh1
Y1JgtI17DswjjLqat0W96S2As8LVoSnFhLL1RMeh0GftNK53IXFQVYqoGJ/ipgs4oFeUDkRzmqtd
KMbYfMZhG6T21K9+TBzoWgK7KFuOZCMor0jRdOgsN4b2JholCDWsfYJoGhYk3fHYJH/xKtLlZLto
U9olT3wbtVUU7snqX9dvmWIR2PyZBSuIil9v1aR9z0jZWr/3KPBIVwruz1jeR7j/wlURkUbHlAx+
m20/AP6KcDGtq/7Ic/C2IXhV+jr1G5KKKjNC9ipPoIC36wd/b5yRh16JQc2EfxPy69n+f47D+l1G
5Syv8ck8dwpISWJaRfPzjJkW0dcxmCCmHGce/M/HScjv8GO1PJORB9a8TGbl+2bSWbWBqJtZGcJI
4xvSK30rE4HWr7B/OMo5uKkGk2Bq/eK4Xc2Ucp2VHdMQIDBfAJ17riwAFMej3NamUpo6MJe8DycO
UF01ofBdproC7vN+43re5yEUFd2GDyfP1f4u5uSMG7urHZT0gkYKNIbYsYkj3t8Sfu/AjbpKP8ND
+u9JrUkYUMPIgeYm4XmeewsjwwPEUgcT+Xwlal9VtNbP9t+pkq1IYNlsZjw3QrpG7aalwBBNru4J
1ZVES0UuwnKTu7+SxSAz1eCtMJ4NhvR1CTtg6CrhQuPgl7YZk1XtWVnxQqXuqWDJO6nCx8882MLh
2/aW/D6LS/Khfkz5teIh+MIjjvI7HDk6sHTSEKPD4N5KeLDbzfUl6zCzsn3sJlH8GZEKm/VL0y/8
vOG88GKw31GnWubAU4HeBts6SoRLTihD3JNa1XcZaBcSiga+m2F39Hi1YOfAOzdKFPnIDoLImH6w
ZkmkUPpVbRpU30GfpbaRgtgKUFO+ywmpG+QC/y3TV9rjWX2GuRjrJQMKiUGwQ4ta3r0gXU5RhOKR
6uzh8rd4qR7Mo6zrMQY24Fm7s/q63kuxiVt3RfLID+hiZiggM55VGvV8shUH7Eg9Dto4kAxoDDfd
bqkh985NlhnbnALMaYWY/IP94zKn4U7XGM4yr4HY8y2y+iqO+bXX+eZHKQFyCe2ACue3HgoUHnV6
9c9qFPaqAa9Lxo100RYgbsodQhgGay31VOZmjlD+COgIwzvAfOjdN3SmX/tJgExWB1ErWJGhgUaX
URx0pgMsBNketUIMy5Ga8fBPqD1IHLOx+LI2SBkNZFCcbKAnWlgKh2OelIUXg17zfCe1k9KDfwD+
tj/jqadxd3k4UUS+C6ONvyP92UAiFXYXCr5mCnkF8CD7/EqMUUyU5xvRjbmurkHgCvKtY2OFOii4
Fdi5RQxVkYv8pxIUTUYt3CA3qCP2QLPq9fX6+tjEJo33wzUtm4mAoz9m2aT+tXf5QXB+YyTjFjRv
vLFiBu66vrpnZcO0Y5J4QkNOHafK9EwMp9gSnTL2PP4WESoXbVYyK5hbhN96lYDItfpVh+5LjtX2
+4xcHHa1zepoyKrVqYo3YCJp1vCd2EbUN9eIOzgE+D6ZuzJXss1jjRqIDnNojl5da+EEzxPrXaN6
hyMJSUyoQM4i9Ocq4tyWHYcjz85hiwHr4HCldjG/lRtOBLtXPqhyIKuy3GlwOkBXDVALhW+HioMO
ZndOClbZ9dUQve5MOfEAWcng4di9XJA0FOgy2lwZz/z2Mw9E6o8TwaaeGn5y0cVs7PFRZH1J1kY1
x+ddg4qaTETQ6j3PgPBvmf26jetH65bkkn9FLrpSMQrtu4YLE8VhQnh8C/FwhHLjF6mK7jJullCM
kE7z8P5Lxw2PF+vMSEAexnfVvFVTlVJy0tF0yM6dHCPLvSqPZnZY/0rEEpq+llEHQUivAbFnda7x
Y/q6mAQK7yFB+KuEd0vkbCmad8pvmDkB6JONXG2h7akHuQiBKrF5lmTvM3xvXEUcTKBk0ZC0IoWa
pvuX3JySif8wUATFc8VC18ByJ/RvT4hsxrlBNekSbmdFWqDKT2kwgKptrYwt7uAAT8kzKmJaURnf
VdGTYzGZrKbajut7utK0TTD74BCjUx2hAYYhLFxjSZkUakARGLRIlTnxVo3+MaxLnluQkkBGpeJD
MTuIUGqZr+11qxIO2ANj1AfORGovioHB7Bo6nCZXzkHkSZzgIFM9MVBJUAEdsTCqZ6Bnx+0yc0YF
PHNACYAgF95JzIh1sPaeUflzMpvtjPcRWuJNHh8DJfyjyxGBQEzy31QzB7xh1oNXmkOXImrqSIDe
iGr54UmgAlcLWTNyX5I5RK+xkPpjXly5EIY/EUADrw4slzwuiyZjQsYWxXlMNiQiu1W2Y5GDnGvP
aTGtIIXkEvvLQ17TJ3bvP7YggXNN/20HNSZSJbvsfP33HloXQRsmM7Mpsni75rFtdDpsXBCFeuwO
UPBkxhPQ8GhgCWDUzm5XZxrQEwMRnYe8jQgKZ73/AWMEBLTGcQBRTGYrCVuYKtBSXmVEpaiyDWvb
sp5/E694s90e0kFH5TLlaFwSPII9HyXtGtq1XjKIuNRNwGS8VRdGcySxqzcgM52L9vRM71RUhN0x
wpZ6S8OLvKkFo6JNUmLi2KJyanpqwX8mpq9LbaYCjFfbRJcSipCC0HY+bPD74tp32FDkCASixWwW
fbZx/JlIAJIEpGddo1mOx8K6rdhrXQqjTJNaJHhJrYz0GaTXNbrab9LPaSuA9fYMnaoB98FyzCxD
YcuBziwLr7KeFfMRt2vNjdB9oCgzJ1AHBeDmR1CfQ+uUfR2o46Ko70mXLQrAJQS2fXgSBBVBHriu
2XJ4RYYjxSfEn/lpTH8GVBZPmw4MqxGFzAk/qruBn+vvFVhDq+ypZ3CMHzHQl1X23BadFgp7VvXd
G2OOCFDgXYbaZYznD+mkPh987Kf/FHFY3J0NK9BQ3Ky3/kBvxO2Mmrlmi6Y6F0jvJ6myKqc/If/O
PQAheGp35a7Wem4u5i4c++ka4hhhPmzLOZgnNbIClV44ExXXfgipcasQkcce9t/dPA1zEx0G+tAd
KpfWfNsSiFd2J/GiRS6V3B2/wSEZ9IdoRWOZ/886WaPjyWoamIKuHUpj8JGWJGkbjXKFZh7FcRIy
n3Bqj2ku4SuDfWQNrQ+ftSg13GioLUadZ1de6uasHB2ENxDWw4XdlBvgFvnuCmZLxP3WC7Pem3yT
JkCAdxqEXgD2g5FisXTPozQVOfaTsLgUtu67uDNJ/3IT9lT4zcNhLuxs381b0mfqsqSsEfJ3r7LM
BiLdRnbMn5AiJIKUvS+Th2rXl1Mi/Crgyzb5L+FMBPiN7ELjfqmgexzfZGS+1CHLOnaB71mg/xv+
cg==
`pragma protect end_protected

