`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ciyztpkfaq9OL9GTxM7O/wR6NGP1yBNzeZYyZ3f7Q1x80+G0WNz+rEx2NRJueJu234VXdcWjqXaN
PaSIYZQqJZhM+DNSQi3n7eB+aHgdfoW5b43IkEsfXARQvqp/2qY8Ba7kWEMxiOtSQ69vRSAqhk/R
+zZByxCRkK4m8rNL2S2NWovGzJ0XAW+aBlWaH92VQVFz2+b9LYmD6j02Ph3jBtAx7G8jUEaQ6T3+
5eKxmHZNr0Wt7tRPQESxWI5Cd1LPkYU1+Nu3lRbFeajY+E1I3KHARMJ39F7wxXPDvwwIzktIPv2y
X0RqVhCVzYdlzupaD9sRLp3ivDDVrNLxGRWQYg==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
EZiS5WkI7f8mcOS5U7TRL1HLK3aGdXf0OiG7RlHXVM0ZE0+C/FiRYcPLp0lKmlbSLT4/vILoFTzR
5NcFWfVWM1miqjYic/ePRH8kDiCdrPaC+YleUN222uVHmniw9E3SlSLRCRG4RTBicawfdQ31cYCM
I+JLk47Nu4iPL74LemfANwgVpNxNC2b89NGN2vz41OfA8Dyt3xW5iFQ0GlcgITydjlbKInMP094E
4nCFB+PsdvNnLTiBsYDRxWHtYwo9dGKIwN10qvmZ0EYcQdL08qZ0mR9ER2a+EgXG9VUL51x9LSuV
1X9hJF0nOGwLDIs2EMXeEaowtpXKEzPicdxxuwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
h6GZuBWjR46vPrAXSs4oIJIBB6mqoF7szL3amRKkZyH0Vz3a7aeG0UzwACSTEfIw337DZx1Q8Fdi
q+XwGvlezg==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bEou5n8u8O6VyDKK0c//Ic6L746i7jYD+hb/Uip3juqNUr3jjSkt1G7MZaQmbHYheg4vDZEne+Ac
4KQWpZkeINmYLJw5AdwLTxt/xYx0vjSCeevD68aQoY2A4Imls8b2PcFkeUcgM++gw+rMrKBbvURQ
Au6zqeNmz66a5h4yAH3KE4PdESzaVJb9R+5zHGB6QgyRBAKm3/oU24VECwinc+d3/zc4XBixVn6L
a2cki1kuXEPERcu1YUyN9BHwWc7NfcZ0FfsMmblXUZUIlzTnFhGCazEgQezsOv4E2fqv3LQsRzbP
CMXdPGMDvBptD8FGQ+cof33w1vGgzD+j4FaYFA==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
axeO+oT1lEEwlH5tTEHrLOEwH+BzlK6Tll0cwN9y0rMdzJiUCQyJsSDd6i6ZCRWIjWEghQANMa+x
0dOwPxMoPIFdzm1GGBcqcJX1cu8C6jPmte45Oepj20XsK/Gy18S+uB/ejw4XMfD2gJ+ACkcPfXHX
GM88FuX0iILs4SVa72AnbCow4He9JUl/lwDqf87rRluL/ufKMlcIAFTGR11brl5D75o3OkQuwcI9
3qfJbkzptOr6Z8TaXlExZxfYICqoqyfVmCXFTb7+QgHkmhOO4TlAgWp085dePg9MpARSLaUByT6Z
Dut8GAp4es58X/nNmlcToBIemTcmlBAXtVJKLA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nk79QyU9zOaPR4Lj2/F2NX64VgNvUlNeqE8v4dsC5y5I90Fasyiwbl7S3OhvB5UPl2AKwVa/ImOb
7PD2Wjm/kI2GrE19cme+RYWj8bQSMJMFzST5doM48CNg7JwK7m6Mwtpn39flxcxBSPsJKoTpwfFb
0QLTb9gAMtN+ZBqxIhI=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
E2NU9iTbSBgWfo2jb15o6QyC3qyj/cnaZON/hv7sH+W3GIjPw2pzaTw4Kq5PIGHUSO2Up/kixJVa
UCbtPgf4bCodHBXL63zp3LPYQ3vKh5/k7xUugMOHq5NG579BlEzBiPENEfBHUtOKNSTTPoun0bBl
NblN7RWQj38SXCnlKqMhMEjfPinbMLwcOGAXPCQnRxlt4RPnuXt40UpYZivqumEzxe+iM7YGVdBa
5a6zh+eAmgKyP6mcebmPpgjeuIg5IKqZ39FUwrhivypbXerNHnLtTCdxJvkwCurG7B4TSLBCoJvm
89UFQTh0rcRjJKrnpCI2zw14wNHXKJfpOCRDtw==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LDHa7nJaJeIS8PUEa9kfmJlo+LK4y9oQ2iat99Si8OQV0Z4r8OJu0Qc66oaPhVcdw5n97E5NJedq
ZtfzsetTUSHWQ1P1cruv527J0oX3AAyNVOpzLk5sOfHyAw0COCy6EItvIOWBdSr2AiEtmczZcUtU
sWO/D1xVMzVnSeU2CLACpQP6tkcQc/Sd1aR7vAuVo7XrgbISljIaJQFxPzHKlpJZ1/prINPCHyuG
VfLWWpqxDT0OTXS5XK2KVt5hPBjS/KS/RT/L6Bju4tXX6Q0m7PV3CdrsPok3GN2YCO8ihGvu6pqU
XsC9QZ/H4gOnFHDgpMY99LYlzAYoLBFoaPj/dA==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
sBog3Mi65T+JQsAl3ryQT1FHV/a5MMb0mfWA/DOX6EpF2UYzyZV7clMtSiEsZAE3vwB4ElhKbFhC
aedhBup4w1hQSZgsiFhFm4/ekFZBmq5FbM4YljBAObaSZPv6sI+rvx3Oknfe2SPbjdcTu4u0OXFe
lI0X4eBuhHNugWHbMKk=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WTlUcdV5+Sw6qYmmuwPwsaC3WQKUa4j+ngQKgULUY1FGDG2yA2v/11v3+4NhE5U9LJ7ZVRrJRgnp
G/NOBVrs0JdkLEOJQPTPGE36rToWBsbay2K4fv3cyMcz2Uan/QvMdDalTtGrYWGP1DeboIIdxeB2
n1YVGWGJIBrW/2Xf8/BxDVnTpvFmdnqmlBCCWVlQ1mAYP1GFkguU3uFsiOl0tqbTvKKURz2FMB7G
CcGHeAEGfl5VTaY4gClYJzv+eAWSlyHh8sQrXX7ALpAhaQodAht8QR6000ghHEUxYpqVOXWNDOa3
fwwwutOubxlpU0sIuU8Q3W3w/w8xCOYpZFjHqA==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56512)
`pragma protect data_block
EfjGODZSgFnmDmJuCHJUSLptjFQNxC4R7CUV7mhPiX+A1b1/i9LZSjcaddXuqfTETDGU3JwEe5FM
zWhhQtiY0O8CR8r2SJLRq4uLEA+69rotuZcxbhT449F9imSglR1F+Ra9CagKLhyLkuOI/0SXPTjT
xpWzLFFkeUiOaxgp0q8qrqsdlOnmmG6UlXQt02Ck/7vXS+dApiy7XDoAFnAa5YfWLIeBiLKW665Y
bRJ2H+rVXLyU9MHW/cpG+RddPLgbxwUGZnI9qZbOwdIVuXC8usQa1XPQWtFFw+08mOHHthMNkT+q
hE5KVfmf1MrMc00H79naTXyEXZYB35ombyTyXdb25nLxSmxIvJNuDvajKUIRkel2GHOL8DEwmpAN
1JzavpkMdUtR4sGmw7tl7+ngb8bYmKZdbH/BvqzBztXgQ0kSl71F9NTpsP9uZ0+oqqt7jWZFcwLC
A25k7rgkYctCgWjQ3QLqVtwdEOMvs0uuR8ZwiSD9NfyNVH7hy5u9mguK1R12716bIctZ2o4UejX6
V6wp+umO5Q5CGLla2xOEnRb3Ipsib68JTPM8BM+Ovk2zilI4heLzDoBMpKu5dvQVdNXyieDWSx+L
c/1WFGCRoBLOQvH09fbLRssYRbYQy5hDCfw28ez2tGxXQwtVH0QTEJen1JMLk6vDKw2pTMkTS5uK
KsKq3dLdina+Ysmwzcr8Oi4sC3gVdXoW7fdTbFEvl2ubmEAK5eaJIO+K1FbEpXIHIqVaUC9KhQxA
WXAb1J0qJ/2a0Hp6zSJEyjIAT9gcccX9K3cAhg44twVPnf8z3HbUpKq6pwDTvLTZ1WloJXGZesHq
Hakx5BXHCYE2D3WnBl3D1zcTXK9qkwsWMmp61Uq7JRwVqBivqoiz0X+ai2nthw3oSBi6i3/fv7Po
vd/M3aENoqW+eQrsxHeyKNm+ecPoHK45xFrs3GH9n1Lg/3C5DnW9zq5tTNoV0vfuZh5Q1o8t3WLd
B303VpyFeAutcE8XPPfMDs3pHX/e43AETuTK+ADAGPY3yQchFE3xEGu4qdVcCCAh4QVsyPeUtwnB
5l8d/M1R5F48gTdhS/1pWMMSP0qPBwoqmk3k3MG6PY3SzkTtwYtk7n753Vit5QpES6m4SgmhI/NW
fGXgybu7VbLc4j5wtBp1hhCEdJZjSS0A0dRfQvVZwXoyidkkIzBQcTv6D968vDJdJXZME1YmRPN0
wzFX20z+9xKu+VbWDoFAlliKi5JgLe/ws7SIfsyVVV4g0KUx8f0uA2SkRMxgiGEYSVNHYCQiepiS
kn/bZmm4Q/f1XPvSOBnPsVt7RYGc3myd/S+fSHsCxc8Ud8M0dAOC68534s3ZZ89TVaRc2MT07AFc
a4B0/yegEx7d5kykwxPCULHifss+VsE7CJC5/NsNdz2flQr2QJ2c+i89AYbXf6nbTANqxIPvRQQd
xasHH2TM1lCvyPLKP+i7885FweDN/Mz01tiWwfvSXm2DEKVn3Jc8t9QFgTu4jKZ2DU/8XR0YFsRE
QkANh9wzRDPF7SHkodHIcIxGhKEQ5ubJsNUKF5zayAgMn7+t5JLyFBia3+B/bpY9R3UeZA8ORLHc
nNlpY36wTJkPF80/yswSNIZoG1HCYY3ZRGbg2rQ6/x0Bdn6vjCPb16ojJ/aisdllqEohviKgrKvz
q6wX3qqtKFhX5qSSB7Xet6t+jE0xKn3YRc0uozCSxaU1WiHWiaweVKT0vVYDCIuuNGChs4k8cEwL
NVk9cvkAXkiyn3ntgInx7qCcee1aMpKl29zmoElbQUxQqflHsMgafNLCGtIGHxBDW6b3ueKn7+lp
WPeHzMtxWUTmDoareiTy7ohAqUD3X5URpIC5IrWkM+Cx2CJVTd4hctOjz3+hcLNQTXi7hPG9LJNe
KNNIf9RWaA0q2v4ufzRE3qd6Ev2wc2eJ9FoXtSyuNr6A6tkznuR4xRpZsy84PLzGAhkIgKfg7K8M
GnMDa0NkLd26yOSU0DP5Spn2RKhfHoChfkVH1D2e82axNZyHf2h/ZDswOHnhwcjpvn+1TzLHikj4
JpT1hSjjJ/xG4c+YlF+ivJURWMvZMM7t/cajnTVdJyK6FZkuo9IpniQWvizNWQgPF9FkztCsJbwv
A0RO8pLR9WONyDzahQPzy/C5jiVgNkY7xlbLq8NoxtpU2c0oj3cv4yDwOPMRzC5EQCmuj3lXBE3z
0qpdDs+oaQweVRHZ55adFx45Bcz85ISt/CVfJBMZ0NzMuSrOEONem4MjU9RCzxTHFAleAtXR4H3r
GlnbYIhoR8X2/2UgpzwqsMroVLduZlLbw1snFwv4wvKLYx0YMjpw5JLdtqLStBHCmXjc5eCVjz14
Co6bU/eY8yo4mA3H7ppeSN4IVyGE9cs2qAuHUAS5ltdthULuQLntIuKFZaiYEG3gwmjoti5lJTJ1
HrUgILox7dOYl9WtEjRT50Bh6ttmMhtAs5oU3vcjBWw8HQEBuIlRWBx6jOBfacOXJt54G2YC7K1R
PRY3gB/Wc8NaEOmGddU816cdHVvf4RQJVbx+CEsJkZ0hR8UYJJQtDLFz/EZM66spKRnVR00iyaLB
8Ltqohk8vdYZeUlkXjG9ao+dvCmtRaxjqu1t0Ni1NlJyWHde6bbOQZaL/U+tN/MtnaNi8CMCJMzG
3ItM5Lg/Rzq+t+84tmqXW5YHI4oaXdm/jrl9n9/wQAL7xDI4+hEIlosbca13XPJ5kEBhPKZuKgdu
icJ57+LKNt4rN8fV/pmn0MvFfaPwypRbxBXiJE778zukMJnR7d9bgRDRW1LeUQNhWHas1gQsMFyh
V4rZAod3Deg83rmMCwBEDG35PZ7V7ijrESvaQAynCi4gWYyv9lcprDyLGvU5EH1QvkMAE8efGwrc
aOcQatct3ee0Wc/OOycMMspQGANX1Adfoijhg9TUuT3ya+J4p7bbW4KJyCEnqk6VV+7NmhTLrrEK
J1Oekvn5qil6JS+kGlOEYv/D1EfSMx2eYazG8k6h1vb1oyNPxl3T3kDIWMFW+pSj4E9sj3Xe0R+O
OhhdNWmbnvcIcV5UKG5odBHIA+Z2lBJtypxS2sFx2NHvuOR8vYAbB4YNKAP90q7G6fCaVM/I5u0/
bCpVJ7C1aoh9b41U+00fNm03LqIxqs+oMgO7fuNY9O6Me4AdFhgrrWTB8LhAfPt7TOe920Bj3A/X
CsQTEpQlsn8XBTyo047L4SbTnb89oVfHIukCf2zzpwEWhAInqV+KoU3341UjzI0EJU7cYu42Y06/
iFK6U0AF7chls2ydkKT17PryX3Cf5A1K8zZMxjySbUnb5ychE4UgfvHHAwjHSesovYt2IhT91lwO
BvxsntL/1UqDcipy5C6oZj3lL+6k1pk9Wk9BnuMU9Ib2Wrv50YDb+G5aSrZA3fiAbWzYF8FDuV1u
2/4E1yD1AYsw6tz5gWZ8uLWlQjvJ+gdvwFkBKN5iMxPSi4hhv9YR6NcZ0HRWW7NVLPS0xE4eZ48S
DLyUgh+lBfzLcCPOvR/Y/Dg6Ngi2Fvaf/N4mWuWikIZBa1zep7P+fQao244L8EKjhPPe6EXfuvTc
Rbf9ZXPVsuMgZW54f4Wzw10Ds5WdEoxEEwhi7wBm+l4XKUfQOfHi3J9QuIsEIM1eM3EYWAcFhpdR
u+llUSlOZqJuOyCpFtXbeUVaFhPG2nDL99hsQy7kc5LT2JqROKufkG4rIkQWJJngP5ZcpLS89pPr
lGLbcMLQ/aKOXTJWagdThVlvU6Dwhn4/RihvVa7psoBWWLKvR7gnb1s+OSiOGo7vokADwIQRsnT0
BY3Jw16LeYK4ZetsY1Ww6wWgBBxs4FmB23+ZC3yeamvaDWuZ/hhZoQffjEe68USAD3pIY7f6LK0e
7K89fZfUijGgdjZCDzcNcKiDNYTPQ/SMvQRy0F97KobNPteW116hWdDaPzqLbZDRuLIPf6tBAifh
YiWLl/jtU+V+0JuSeotivSYvftBoYMzVCKTAA9OTuXod0WtWyaRQhV8sO5u7nczcqcOUQ77K3lGT
wCWYAdDGpQzFCi9rXJ275Uu6hOULu7VMTWsVB76n7+qemNnNMR7gK/cOaNWwNi7KKTw2+UibiLXy
66laVwJMkOz9JJF7TcO2WPBXiiHX9Bfw3apcTjimB41rmxVy/jSfr2C+AhT3C4F2RihUtFRKuk5i
c8JM9jLuFtoc01cEJq1QFQ4j/q7Vepg2Cx1LHt6lj1nltji833DrVHmR2SLH1TiRoDznrfkg5nHR
yrvmxsrVXEOXSrXCJSnxN+cZUkoP0jOX5YP7G9iQg3M2zQd+BuUTyKJ2KP2QKti558Pu6FRlk+Se
1vfwBGO/QDgATREdSLnCqDe0ej5WTqY+etrCxKMQMeyGXauFylX8YbPe1CXo9mq01+JXr6torLLG
ErKbLqh67r/VTR1JoRPr9pn8X8BsvkIMMsDfWjCZc3UG6PYehRXz28PTMDwcEN61eOFgzAtL64sb
j8i0RG+JOfTvX+4LqvkGftSx6sj9KL5B4WsAauqFqi0lfSphLcLOcpkwQyGG0uGoHTEVUfatWCrt
AaTGYDUm+EBgzR7b9DmR2Yk55mrajioMyJlFxKhVZN2WDQ+PLxt8WgY3C/18filcIJ3Q92p/fns+
V3YHK1lELKkFY61Jfc4p3yfRKdpzPehvKn/DpY8HYS7Aj8ZJdHjcFlpOONSn2Wx80Iv1QX6gZfgk
KgCM1FF3emVbTr4Sa3g+b+QSdhCef2xr9TtDN1TYq6n7ErGAQFFmmCOMuHTlDc8EUPBlAWRSYG1E
556j3E167Jr6V2tQzN5/nsC3t5//rgd835mMBbKEXb9VEHgtEn/5NTBLQqpyYbYQ8K620HKkiBdl
izNVRKmU1puZ9UqedNrWwEDU6Ly8MCa9adwbeIIn4pCqLPmqJksyzmkz0/ApGQgrho/SrgkDE3vW
TEMHXX5A/wuaFqx/ro/4NQW7n3NGZWHTYqh6thNY/MfSfTaoq/VvJT9m7suwZxBR4lR8dfhdOSFx
ye0Kd6/lZz8YJAXBvRFcwBrcKPQcMPib1kstZun5lBa3sOcwtMzJ+DK6j7pllsCSQHTOoIiE/arv
spDXkTD7qcBFEj0WNNVUcZ3IoHm/bk7zVmxCtnpgDyXsBwG8lk2Wb2u8oMwjz1yNoQRbPNFkNGFm
3P7k7j/rsdRpFYe8MaiiM17ZjZJv/WHRlsLkwLPfS3UtymGu8X83z0w49i2eeZ70vlUnS3ael2dW
k4wwMfRIHucF2FILgeYZQrHYws0QLKdgxYDIP+c1CAIzCAaF1ziBoI4EgA8Mu4Xb1T1I0bS3UmGD
f9PIsc+C5CHGZkceWjuSuz5Yq4uypnRDWEqOe6zPQt846Hs0gEQWufsEXj+WSe7KDEgKyYloslDF
BluY18wJO3g88N7h/EHHKse3Xg1iI+9ZwuvMfq0Q88wjvAb+w+bGfBDR0D19e8WntFjB703IKQoW
IVOWwgThVdw7cAbUqdpBnIDHWPMxPRtNiiHY2WcTdh2pqn8PQNE9bgUwZxyVfhwmwlknPxbqI5Yz
tIsw78PtciRUcBVd3p1/pR6ivrLIBnoaw+oEcqmXWeRwIkSQYOyr4hmFEUu82frhGywIjjviDqyv
lgcxnhmU/pnbX5w+G+3tWK7P9rKfcSGnnxPB/RzlHlMsHbaxCmC3NOiCaYEPnwW/fBIqbehRhpnk
1kIGFZmxvv3vYFkVpPYwI1tCUQUTnIehq4F4tcg4caAzzA7ryvZ6n9AXmbtb5TozqVcfclKNtPpV
bx1DD/6r87FPybNeW3pHDVfDyc8qA8HgHsIYe1R7TlGd1sIocIw5YBQ6nTVFhWCsapm8mc051aic
eetcfFfPaBlEc4rSOGH403xMPcSiljGbaC4Z013VXezs64h0C7onpPUMTkJpgrz5mc32vDLy1ZWF
/Z9l1iUsfwTlbq/YdYPOal6caAvhuLX6L2nU6vvcbwELmbvso0uur/jiUywTPm+51uSrOYyEP7RJ
vTcAKC3o7vGKJQ1oWqL94bL8N/Kb7+INIXn8EnBcUMEceo4Lg4v4mbQ8mLHJXJP+E5DxE5jjVDt6
SBFoqVUeezzYdCGA3T+PSJ8dClTyog1TfAJ+UMr08fd97KlNVUX2wTyf1/CEGwCYcMhGX5yqfYfe
Esm0dbEuhfXIOmnzV7hSOWKfQ+TslODzOwo26vTZt+QHFplm8RLwA/l3qu1PeaHWt8fYu4949uFP
kOZUvkNuGUSjFD7V+B0e++EY8qQLYU5RgK4wumEtLPz2r5NshVGTrA1YlLiSITHpr9As+HaJaJkD
HC70bZ4qRTBsDz6QCDpRZTB+gbcIoRDw7PN4KzmDS6PiEJfC8aBAhEdXeQ1iUu7Axn7B//eKBtKM
1MOFz7fuZSe+zvUHMdf0jOUOU3GH6FQeWW8tMxVRDHvWF4lY1syWu06AvAciq4pPFeuG8P8pl+ke
APQetatGB18reEKUFS454/68yGxaPU4ojRFs0hrF/V2Ej2RzSLhklYzhsOkyrOoT8ZIGZsVkqHmM
m91uKp63abyzzqMZWSwNTJuAVG4sirtv5dCxFh6JHB4Q9HWUawcjvyMWHt15Fc0GGNVa6CtEi5+W
UGzAznEQ2orUwCaRDf/IM+3EVeKun+YkurjgNHjWbr36k5Wsl1AtISEKIYgGP2Z1hipIM19WooEb
BKDHE1odLp+UYZhonuEgaM2eADNgzLVNMpq5vdkFNnUhgmmnCjXRL7ox7fhAKBAI9vXcdGYTB75I
dWP4E4o/nLEOSjf6izilI9TeiDkH17CMDJs2Ba2ITSB62QqOjaPvIXIcazLhYvyfDz/F78tvqtHM
uXFENhnkcbmE4c/IKihKUU8KuvjFSkxoZ/qI+SdrFXwFeiDVBbHcuTQi1/OKnicpBaCWKs/ID6eA
RfLTXzdgc2UKPUOTiJuDMDNqsSFECO7MPRuEuc5mR33cakkY3u2NOYlPhS7WZyPx2cNiGSoxh1nX
1YDoL3BKLmpCIwnVti7n+BhLqFbpITAQOZ3LZczZaz7nvt9JCKtP61fEUtvFOJ9WtdKmvlcbRWgL
yXAac0NjjVyS2MJhxKlQL5A6x+2SYzreig25ojx5P2YD4IwS2OkQ2HextguGLgpnVq/8dDysYYnP
ypV7CqvE53BNQyzfnZ5zaoK5Hl6UWg6JZa2mXP10G/w0TkXIiQmvzFL5O/E9dr9/mckLFt9jPQqO
1HiCbk8yV44IENfO6mXBMKqrRye9eusbTOSIgm7CoBFH8Y9RXcb1IMuQU0jBbvLbwyqJ04edYn25
P5VZBU4s77IZCCADXSHCzRUVutyrfZXaFd3R+4IXgPvLec3TwEzamZLWTcuudCL2LkpPJknVRrsn
rFMthiVTqMqfPIi1/9+t111rkjYcMgylP76onRzIXcQwsBiXUivTiDd9pwzWMXhPIy1QFipvdrf6
zaZQiael0iFWN8OH/gt/55lrjHSJGS8sYShcldkAEfAqwzDTn/1KRAkrOmw2LdfST1B7lzY1ZHlL
TUgYvovwwrzKtrifGptj+ikICf2aEYUj+7tR3mWsvsIMJBOS8G6puHSRaVJs44zQbz+b8vGAoHDG
FqAaFOm1I3HJzaMoyq0MKny8N/QmKaX9FBM0aGEC2n50Y91iswy+CENyH5zUObSL1uxJt8Ds2mod
pEVCItZ1F8qy1Vm/veoc5m76bVawFzb5aRfNcp2EeDAakvcMcKI7hzPLwRogDkrCcWp/Wh0zVZCD
3j5p4czDONl9qAWP4NOqS/u4DwHwIyQxuOUwEbo6Vqpm80rRs0apQqLuB57XALnkG8n/RLzkVacr
cDkknR19eUkqLpJWnvLFLQeNxJdKrt6LMDGlBXqe0aWCciOWPaRSAJTHSLppg1/9hXTQXny6iB1Q
1UjTd+wiZsEv+kLxT/0BiSOnWZwFtbpHQkBrBnrqeDucu5QVbakitTyp/ow0FfpCue04bCJuF1W2
WpzSbcG162BnVtDrpjs7Q+3CEs0mQTYSev9pDy82OrnU+aBgA8anU48mE3U87a0OFohpSp/tM2rF
mKiSODvu5d0PFgaVNjFrSVNs6edeRr0ZwXWSWzyDtJ+/mW6HHZcsOxrLa3I8SUvyuhWC4ZXPcZAc
ZGU7cYqauDQiSHyalGsObBYguixTbS3mfgkApGXwSZ/FkN2KvSod9bybrpmdk4ZzFgpjI7NqQwXG
7z7nHFJ5GXuvuc5rvhsaMvTYHMRtTPqKKM7Ei5GuP/ZvHpJusw+VfzULdt/ftMDJIFoZs6PCvRr8
KUtZaCPceDqsYqgOQbiJQbQdU5ImTuUA3TyCWeLo49PM6ZKXzbbcDkUCjv13lTiOG5UoOqD8fOEC
zompELbHgl5F+dTqPbNmK2+uvUuiF14JaOKGZz7hwSUifNs9BMObU4f9L/EonZJHtao5Hislq4rP
X9mE8nMz1Nv+5KB0xoL4y3bUoEmlGputUJ3yZEc1nNy7+LHmQbcOMv9yLB/kBMM1OFsyj0AATO5d
gaW7Z9ofpOMKapoCKMRz4c5h3oK6gZiiszoCqfVboJYicv0gOzQhXMcralQtWrTscMhV4RBI+Slz
zBpxwditmc3lcANzm5k4aUfTuouQILuuVjUNhHuQY+yT+QQcICaOGZJfVUeRHb8JNgXZ1hg4o86c
6PUh9tr1hlSOFWjnhYugkHq5qtK9Bwbaa2OESuxUZ+UKnsdLacMNRAFVLwkH3TbcP6GW0qzOL9sx
j9xPX2a/saFaeb2VIBhjpvk60GGHFCrOxE6dV6BMT/O5GVCUJGHxagzZvvB6BKSgQBiQEKUfQ62s
A4dG5wePCVIZtxPGQxrjqXFC73M5FvIWuPpXwss/G8vklZmPA5avxg89OpXXCHSU7EPcz+bTXl6S
NooaU59ghqvCkDym4jH/oib2Ga4tJzOpCr4/doElpPCE0CRU0YuEw9cs0TSRFmLxT2quZUz1PpyY
m/r9XxN0aGBOOByNlyqMpvhFI7+VVOWLZv48GFVSysy/DaLw1+ZDaEQY5le8/q4liPOORE07XMS5
jb2SW6eGz8uY9d5NRMfkBHjfJSiBKWm/bOfhU8ktiZ1VKre25e0DEiKBrazNuWyeLm/jxOb2Fna/
Dx+9B/WGy0LaTgzM4SBmO9e0MMOvJ1Rybq3v1zrD53PAuhg0G7BCW3uhq3LOi1kvCSESp80U4pZQ
gPoU6NHElsBcjn/rULfFWjIZUSgRGYxLDeq0Qia+R25ceUwH0IZbPxCUCTEuZ+4dvSJKouMzBCEj
8kPQ3XFr0GFczPiO35zoi6FGKvGbzx99pa+eejHNCEnQLNbJkAsTkMlpUAYeRzGwEvqFXxkGeVy+
SRt00jD96gQCSi69/RtVhxnI+Y7a5d+t5VB1Yi6tNROdUFWuwBm9Pd6n3ERhXa+UJ926m8H3MtRF
aDdWmWWyN8yOZhh2kTaDlKCb9ofy6h+CQPrgl7LNcUpPa5POtcK7+YD8DaEtmra9vAay1IH3qlss
OXoCbj+I/ojjkebBc8Xs7Kzl9qmpCEyKFV2yx9ryFhceiwvY+URIRa+bUJfbbQFawyh9lBGeGGRs
abrFMTKO3GJFtXm22KSOFjf+2O+Cm2tYHm4R8ZYkodNxdoQYoPEa1/1Oax9pBLxbdztzT9CJm29v
/PP15Csd52UAvx/oZSWt2JzJQUw0IQIokwjlVqbwAlbzAJyASWIptbAsL51WioZH3QJt/mFJoyco
nsd+etOR3P9CuIScYLfkssU2Xg0y0uDMDlQW6dszy2MsXKNNjMmy711/r05gwgXpK9bV1uiEcXUc
YX9osS4gxS02extbewj/ilrcjlGH2NbOo2GBHtGuvX2gAYZiGCo8U3Heaj50fbQbYMwapl0ol8X6
w/HAWUENP+pHul9ouO3Uztonvl5FRqTUhnLWcpnFJ9hvXSTmfyi5Pi0E3rHW+a2Io60hyL1ZybJR
zMkAWY8VbnfmaA09Y8GG748I7asJjO/frM+pzrTIR2tfSD5SIoMQpmFW3ZI388neJL4c4mBBTVyv
2ldT8HSEMTCMj41TYv3iCPwuvF+NIRcjO05+sEE0E2/sqmXy+8kR0eWNVKvmdjjqAJhDfZ6SkLWp
A6M9mAJ29qqn1TsqyNF2ysglTTXGzcSju7oCw5GD65DnB+KBGbcU8pcdUp3Q6wbOcjFVZ/15LDR1
f5sh/0W0BucJdMkoYvUpy9S1v4DlBBO+8EsUoLaoRK75bbYOQoEI4Xn8FasLUG0FLztw5vt7OFKk
+8taOdXTsUMhVbdoeUlRZ583O/2VbTYA+ZcW2nyfEI3l9d2gTc/989QlZGCMn0f43TxWEpqKOllZ
cC4M+s5pSPNAzgy86KbktYl+vcjTmrc27Y/Trk7oaLSz4d58Ozt6VMEaarhpiL+n2njPuzImzyy3
U+3EpXDeU1mwqv7f/hFDoD9CdhPU7v8M92HSrp8MKTf/SaQTfDQA6pPzuI+fPzYaWdnkZhWav3IH
TlfYvzXQ25Zw/2OD0liG8pxvn8bf2MfFkYhD+n7nhVntpMUq7JqPd0Wf4dMao55yZIbkekTTppaz
OBu1iHSnAjtvtpk+YjLS3r3L3Q4kfYwG86qFHw6ZI+4EQHvti94ApXNT3kjGLzdKZFH1C6ZcKDIr
gsxAts3BnPwiv8F++J4KVFEggYeEybNxsvbQGyZJbgWtyGCHbfZ5iJor3ZEtebyjnhhHl8wUcp/C
x6tQS7gAvS7sip09nm8KXWksiojXSauhjeLI5dzRiVAlTTyYPMcyM/2+jI9PRK/I3ioQce5X6bI2
w/QqgGddYFZGKA6gCaXO1LjQdjBkEr2xyV7j2jNJqrSsa1VwbiQL/BNOVlJ8PrU+EBRnVGw+Cc3v
UtcB/nI1odbP6OzgOFIcYgUtG8D8YsmhDEQdQOlaW0xNecWh2bPeVbuqSmqL/5ymom8CobMiqbta
xgWk2lm1UNnb95j0jHTYf8lgM/9iLDVQxYe4P/Dpb2guItnDrUiR80TDR/C5PIxzBzTh569evkmw
i2+QWoAQUMdRPNYWtoGamMrt+WTyXNxjPPxk+jsZg9bvNGuQDdhUz+7xRG2UjuJMTrcOFxcQmr5u
5/C1Gal3wzZ+KUMdUQK1ohCnHzLycjWgH74EOODm/g1CwkFWvbVllPqkYFpTa/HfSl7LeBKOE8sA
kY2W2dRiDu21x1ANPiR1tHLcI2McCVTauKFs4xLUZXOopFZXze7aHY8svfr8Tb8pq0L1HQRbg7qd
waXoufLloOFicBQoFvAVkdyRmUE41Q6BrnHOYoJYGETloW6caWdaMQQfD5actUKR0gJDJ5UQk5kU
F3sVGpJXpByATvrbgjGszKitzRmkjxJnlAmAZunHHLpmqyIJD8u2zJLkNCHqFPpiHXS93wyZAHAR
0++5pcOIoXCrIjNmxhPwp05Odi3yBLiluNd+qxenKeHP3N5lTguyZzMPKOgKfv30BMgn6typAMMc
O/hZzBQu9Id8SDPXAQdKrtHYN3iW0f+/xeRXKpvcmDab54UFlwfU+i1xeRinOsoyOGUhu2zz4ppw
YDUQ0TMZeT6S/oqzYhMTJ1yNnRfycD94KpPcDfxkBwIB8u7S341ByacFPtg8DHsTpkkO09ts6AQb
kezmLNJr1NxGWc8mF75hnePw00ougipBtiAZWdcg/uEALkze1XTyJLUF+qSEb8X/z424Cm7Abuln
sci4F+t4s9yvieQ3+9M07PzKNRVEONLtIh6vOJ4JhgzJS94uRR8L7NdLDU13UYYID038NgsuCXAZ
Ffv1gwPWUczechBM9Y0PPyWEWKHrzBB3onmcTG8rF/DzCB5PtFbhX7pOde3cAHchPNcxcpilE84X
sU8Yk9LZwNCB5+7vfl0FiwkbMPMDD6Js2NPzeyHkBsvtyv3PX6R50gfcKHACm1duHSFt1pk5/TNh
Z4kzHNjqwgC/KVL+O1h5nDRmZVRsp22cyiYwIWfNVngQvRZF6jFpUzTYYAmavOyinF00ToEwknLc
fEVqcUbj1LCKbxiwkY7tTH6320ugbPEN0uEGOX6JYMx8WuxI9vkB94jYaxk0ymMLNDfxnRExoUC8
dkThwzh1CQZ4lhyiDpvdUQuj0SAgf6OEukIALmTLoj1fzxOHQSDHyf9sM3PxHhVZic29udego6VF
U8HO60+57A0nSVVDSMZU+jGKXXhpr0WgscomuZ8hmZjt5CQ+0ASg5TpyNFbWRkLoBhev8dw2cDBl
WKa/XDTHg7Y+HsnlUDDfxbsyhbomVLrxGd10FJiA0stvJKtqepNKgRf611iqhfahiOvp+5+1TiD4
PMLVsRWbLb2OurJGxIaCpWCPm8iEwMZetu9Xp2xaoEVKJFxB2H6Y6lOkoeZ9SNCsByRGjD9/vyb2
bPiMAKhyr/MO0P75XPBH5SHgNxPkhHKijjXP86PinBO1dkhKqvZutPh+cvpJKe0otfAJoY5exk36
LRqRYiqR9RcVgZ0XeJyQgp8B+R5WUcu4LYBqtcmrNQchrnFW3LmUPw28vXty7qSxd2FPngJ6jwSg
1wJGaKBmihW3XfHex2ewYNZpln5i8cffnV/qOZBXBYo8vFBWWk64ul+6wdRF0D7E0c08AJ2mZdaX
Ye/r5inqWGDVMr4t6St9Ub0eih4Ryt1md3bJ+flYAedW0b/kJzR100Ufsk1KS9/3ZFtE2gJyFpm+
AvDApoqDocX1qPGgVR+1vJofefTvNfn6RSHEEXU6dc/UH8jshx7XlCLpF673wzxjBpTxF1n5+ogE
e4clBoRkOwJYKouTZZj27iW5UL4Z5GU+s4JkktwPYftIzJadZzgTzvHbvCau0XMtT5Mu9Oms+6RZ
sTDjIVNt2HLkZXdpR/vY/YRM1XWt0968kZIoZrtV4Vy4OfplQJc3KOOya+gWapG3G1x38W6EFltY
gYkcdtGq/lJ7KTMuXBe00AscaS272PldfPgxq5Ihy7RMD0cg+WAkE7TLOHsGiFgCrT9DDTa6iJKd
KdRbddI7SNIJtFeLx7o5zd4lXuAlwyMSAMRG0HlN+HxV3++D+8br3kpswhWfvUqkLu4uvXOu/Z7I
lp/kg+J75NP/0MGBNfMWFDk3PSYjejJOHNuLnIRSEjmbBWkMjEcxwOlZeosuST+SGktpFae1rD9g
Nc0cdAYJ8t9XEzeY00egfqc34ONZMJnfwe2apePjx5jDtbo3AC3mP8rRnwaniuKdbjv3wJiXgif4
umJ7/dHQ7HApMHOV2qBPkkIH403pCOYLnpzySMPK7n6vTikU5fiuKywRDIVAKDmaBiOF7RALpnCb
/QRsZ3HjcgzJipjBkhORgBFnWngQvb21H1y51c8n05Ld/MWTGTFfYE2X0jI6SP0Fhk4uFCrGFDTF
H4a96dal1kdhaKs1HuBCfvZc7YDiIjlKuuoDUfoZe7WSVOvo+K9nB/+OU045mZN681UNBi0sLQ8L
jqwdAjIcTQIuqMDAbBW8SeGCrnBxN9JM1T+nGivefbZn8DkQ6YQo/txejpiJ4oArcflPDOHXKjHm
V2sZeLaTTmVW+nXY9GeBY4T5H/mVVMalcunq2IzoemxRlLvVyUkJZJyY3dHNHE6xnIy+FvFWNnNt
ktoBCZXWjlDpW6NhvJkpIe8I3vEBA9r/EjyP/Xw6RdcGkOBMHZGMcmgPC1Y4jlk3hgZe/90ejJS4
qdxUxgAiEvzYXUPpXIQ8hDlz15bRmknIhmkHL6KYQxfwuyXgrbZjRGLpaSNY8dQDA6iwfliatG9N
Ldr3VBHBj/CJ3wC+q96fNE0pRm+ZcU47CVoHrYtZ5DfbT9IFmUAYUpGAFN6nOnip580z0R4QBnPf
Ln/QGFvikFo3mkndXC7l2nb+VWOaku+Y7VfbrFYOQeqAAy6T1YL9jtqP68Jnsvpb/742bEC9R6YA
zRpNf9gJa1uar8RAKfLHw8xf0BknHlLI8ZrfX4Mi7fkpKWe9DnMQyp5BPQaezPsxb/f4Vai22ARv
/PQXAVBrEu0Ytbxl5MhmLjsquMgRXOg/Lc4gWUDEPGr4zGBqV/msSqM7DHLhLDc3F3OtzYiAHRT5
al2lwCfogbKbqdrZBEXMifJzzS/PmeXSXlqbVNGYjDim2lqLXAXsv2QfKS3uRORLh4qMWkSANUa8
DOxV3k4jZClVLhYNa8DDjkYjcBh0Ih7ojW/vz3ucSzrlMlqoX9eX7/CGve3sbjA1LStxOu3dmc4G
eTxAF6GBcINIPqjrHCGRUD+aP4Z8AlMyeDgUkpPu1NmJBCc1tEXgzmAOI9jxw2nArrYu2RqA4Dgh
AAfo35TFC3C+HaXxJoUJRln5z5fcUFKj1wWjtVbVE+K7Hwd4xllDV5eh/LwOdBtsr7tqVzVjmccH
rdxQNYczOxNjCKFsRalsetWKyoP6NznkrC1V87aHKXesILS/PMohszE6PKC6lNAfNIdxUqDMisaU
rBG6Gnw+MB/1zIunJDbyGerqXgSC5+1/fcHb6CUB8Dn0/DRhOehNtE+aaVJt2GXpHKiAYc1Qktpi
UeqefkbBV7giZvp7FM8yZ535CnOqHBeY/TUyEOgWAGa9NE2gY1PBzTQbQKNj1JuBIPc9IoljVK+Z
y5QSYyJdvyAXkK4Oy4IEU/U+DN9tNvsGLtyyOBe3VoPg+yFoMtr9VW4tAoX/Sr1LONo7wMhABG0l
fmdF8Fl1BwAWNLpWWCGdWURUBT7RQWiRtVK//t5gu+mRKb1eykuhYYzx5jOeHQFmSWD7Ax/FS9JZ
3bhVAFtLMj12/vratV/Oztv6P8+BlTYLyXpVwUMMX8Ahi4LBPUsxm0/lVy1qJ9Q0x5uc2pDznhb8
Y0U7n/f0xt+LGiYoSY3V9QbhW1ZKdwhDboeh12o5FkffhfnT/ERJ6H90YyCAFQTKNniF7x06x73o
wp1kPAW23xlotR6zOMr3EWlb1lL+oAjyBK+dQS6QASPbZIS49L/ObCzAX+vFE4ihDlvuYiuLvL63
BCbUJdu9R297i1N9s5V4OzFq61XbtP73HzFAToSOl2eYvMGIAoLSVkY19yZ5HdD9IkrT6o+i2M8w
kpu31SwfEaE7uLaaz7VkPspjybHsZm+L4HrYaf2rFFYVYqaGKJr9+E1i0GSi8G1IrQdoUonefb9y
eGmhHbQ3dO2txwD3i5lNPVBwgLPI+0mkhADpFzYrXRwmrId7+XOC7go2kJWetIwdFR71pZmoLxTT
JxdsudWbtGgHT9r6tVuIfbx5yvg0MBok6Veb9zpo5SI4okZR7oDFwxmmtL+2S3Yjb4JK+62XgpOr
f/+E+gtBsbz1TcFqcEIn+KxvfMrqeHdwGX85A/ghxX2m4yZATYZpTg/e7KRsokpOzdFHthDUBNCC
xKCBSzxwiHAoik+ziwpo1boKIfH0lIWdbLCYkgyn+FrCiJOhKv88Yh1uDQ55c8jQZ6RYdctmztAO
SDURKnjKbFqTe7+GNiWuCwdZM3N4BPDnMppxziDkdWLAm1zVIQslzp9YJXHl4j8MuC0SIoobJzTP
sWQ4dRNIf1HLTduGEGQLsRuH6lF9LaVd5b/6hgitv4xx+e6btk/k+WI8N8JdrQ+M2t3uZPK/bTKo
OeAAni8yuSY1vPqL6ZaEz+PpVL5symUi3SZpf6/54PEboO7ckxQrAlD1u2S8vp0AXZvXYX1w7G4O
1lxcnnBZeAQGEbXjES77+x9g0duVYMHgmxz/YSbMN6E3X0Gkpe3BX/EqGdvX+UfjBIm9+8P/fjIo
Qrh4DfN2B8seAVM4vKv/i3zsDk7xBti9V/y5fXne+t7/VUFpoBNOSQPwsa4t8e7wR1JoJlZ0mzJP
UIU4dCm6+lWTDluKBcGy+SA1gLFdS2J+fgsTo9ghIZ7j7ZyMqYPPjZM18p/YI0NjZtZT0oRBCmH/
zmBF0p/iSGdl1Buq4IhykL+Qgw1fxwSpJaMB/r0KoiDCANlhrGs8vealNf2fcGfve6jVOYSSOcFz
wFVvcoT6WshUXurCu0Lt8KOmlksU8DJDOSb2JMgeSh2wZ3xpcTWI/3AE2lorMPfqiI4n89CM/TMZ
90NX+09UfmYmQRDqJTxWNoAOiOHUy7LDkB3tvU4/+FJJBrAMJZdSLEU87YCq1ceM5j7Z2RaUBTAf
9EFQzXTzGmWL0O/qEzFN57MyXnFavwfOn9cciXqH0WolXW2Gc88E3oFrafQQZVW2GctIEDaK5q+J
V160zJWbkru+igM6deXfLEeGSisRE+1sF31dUGDjFT77yZl6JdbhLdPpVPDyzvmLPgaNkca/g17v
5oAQWw2doIVNPuR9QCmANPMWbyKtwWb9AFTxTlaJ7h7Fcaf/VdOEluYLXzr5ptdn0s03G2kUvvc4
yonLGnxzeBOO0qisp74QSjPLHiGYlEAhlGe1QP/S6RFUTnRvLpcaRga8yoQbPoIbtv+55pxD51Mi
0A6pnIwitcKW1ihzCdgdrvfs+X74z5Yr1+dUV0qmcko8lYzvDm5l6hvbVIhVMJA9m4tmSrQmcnx6
qE0ntc3/f5/gG3HZCWjHmtk7cuZuapctzTdlBhaCy4yIZOfDRLjn0NUOuCQQDQrBASnSwNt5wmy6
j55jpZGlAG3XJU8029ZNkcw6qefDOUQvciXShtgYoZ+aZPws5gH477nMoIVKg2ixncTLT6G1c6/+
/pm7zMnv0aAezmSeTlwZsCSQncqEnbFI8fXos/9CazWowyk/LXayVxC1suoAfCLmlnQG3xEEHQ3h
k3sm7hJdeVnE3+DLA0K9u8E4MYowQ4h06h+Ri8YKb4wlPXsvEYPxUIeZUNOytGowfKEaYWn3dZ2F
rgpq1f6qefD0n4+qyp7dNfFNI/0dou+w88CUzfghZ4vJ6ntfsPe7K+HvF1lLTZANcHpLhJiHM8Bw
o7/kQ4wNB+Z3iD1KBV2EDcY1whjBPhf/Qpk0Wgd6EnpKp/6j4wtRtVPT84IN5oz5F5sQ2B/qnhX+
VXlShfDzlEfiPQ1M15yoq0qH2h916SszazNEYDNWSx7IEZqRHBOFuXU9XUNGAAydi0mx2y6fPYRo
0crnoqSOUBtIXcl0jcPrCG1i5nDGoa5rx/Pnr+pT/S8PRsY67cG3WAjTt+QEVPIvYI1KErd3+YVk
3suBqlRbGyN8TCu0lt4CMzJUJZGkWvsawNoc5/05MgcdGE6VRnwZHjuFsQ24+NdKq+JBlGsYk7qq
pHcRhyovrbVpvgh+2ueU5j7A0vic7ngyD7uI3zk0TJdkeS3v31i8K01DhG7NIsDgncfVHYTaAD/Z
y+MUcyRE4R6j6xNSbCXL3mTxs03TksMlkX7PiP8Qw4kSaPAroqT94/nBCn1GN/Pk7iL/WFlklPrg
pg5RFIyNPfSJ9j5lZuzkKdGc8DDf0QRI6pPdsg9DYC5m6Wuz6ffd+4Ysw7obgr15Tj49Vpi2Q0AH
IDk7IhxI88Cluc+F5TXkHhPMbJwyLcoN9NO/DMN1YJSkK8Qd1sRi4bA9/9MO9uEB3cRUnoQ19yJA
R+DVtvVjBHK8jhbBv0rQ7ACLexFKMWuCsyz6QOzKbSA7Dm52S2GRFuVXlFARe5j3O+h8kMsAddUX
i73Htjm+WnWsG62nKV49JRMg5ORnmfiEhSAqpirIK6MyIUjm+cx9SmuIwhDYc4nZXKFYs5XSo/LY
5M+lorYb7l/D8a79tIV3t8VaB63HPsjm/zOTHtbPZlHarvFfhshdaHRMrDejfCwTw3UjnlWPCilK
nGQIAW5szmawfomAZbhAMnxrJVt8JfhqpE1A1j6OT8yNQnTIzJ9ITd1vg0xFAuMXLVWLn2SZPnW1
2aTNHRHvAxtbGnGSI11BgNvJKTMenRxM1u5F2xI+k5wq13rs9MDB8RQoSf73qHOIpZOWY/Zk+TDb
ldkDkyp07MboXo6Yo1vnNL7aUXPkPlSUaptzmM/YEN2WbM++ftfmOgJlhDpgloTSmxyI0t0qkRuR
B6VDpHf0dXTZgWeJizrn8Gc/tfMrs7Tf0Ne6dNpDQrCuHtjuqalqZspamb2l/qz+yc+Numo3+TMT
lg8RUhFuGYb7nmV5o+aLNpkZh/MIWRwuJwWwnBFuhM7JX4HheOW8KHLJOxE09j3iWeCe6V/G3Q33
6fqXrPbUaN9kc47ym1rORVRl+Hh5sBd1XcDtHJK7ZqnmbIY3dZRDE6DETZGPMeyKMTs4xHjsPejD
m034uDRZzEoKyKXd3cPC9HhPJQpfrMgpSfU2c/ejFwmSvgJxeW7pXKIJfXfPgzONNbD+CH9XUBZT
HFiNCfohKyVDc5PfVD4C4YuhpdvdqVzL4QsCRWKC/M2afuyzho6rYj9ln8CEDwNqI0YGJckQwkUW
mQqEeNH7Zp5j5QVATCKKd1U2iKwLNzTL92HMMrk7rr/zhVSW35lB5C7daoBcupR4E9eZ7JE4m0RH
F37IJvnHiwAmUpCAOah2+2jpJAQxyfD+/wJTmfPdn3L/7mZX71qTtXVokHqNjFR2CuvxbpHaRMwV
LPXy2ch98md1l1RlnvRe22oU5CJNSAXc1a1RoO9PpwMtKiJkjaoAwmxfxpDUacplEnKH2AUO8Sms
EbEP/mRA0e5mh3cB5wa71xDoA70OrtBMR2AWVfiAZwi7n1j8sqSOWBfnG4C5lNSDUzTFeSpoabSB
FYyMvtYg34wWndxN9y67iO/u4Mo2ZVGPEtZIpISh01CzzBLRqIfbCsh9YptWpP5Fg/lyLfV0Mnkb
HG+mIBMswYBzL0fBhZsTd0ElictKtH6Ykl/am+2fQL52DFiM3PNoXdtjLdsF5r6nSBUSZOB0B1co
uXlZYvFqfMiM5R8cwWyIlLN6arsFyrl7C66bu9FN8CO/Ct1GZXIM2yNqo+xMfl4AWywgXS2IIuzW
yUUuBIkUNi3hPO+vC6Bt6X3+Xay9zJQvOF/1qf+gB9mf4KaBZ5U0W0WuozCGEAHphekO9FyFUsuS
igaTcRndVcc2hVjAAqiifK5LJFl5vsy7OG7MA0dYYugMpIYLay2rQfzYK7QvY7vapsaj1aZZd+F4
EZtZpUkBOJAIbCAcKVvA7XvoQhKisxeGnCVcX/BcWC1iVPaYKJdg387E2ILNBkiSTX8t9pmvC6Yz
eq9FpzwU0yWgJzd9JC83l6cahW7UlEZFA24kt+W2YFB8kXtviuMK0w5ipy94ElMBTti9K0EDQkdN
3Dc+W9edviuqoSDQZhtepF62XmyXX6sV8anmeZzmlF0Sp9TdlQBFW8nsaa95IZv67PfonwKkjJ5x
lWoAAttZ4SKb9IpNqVNayxdn946C6ZN9flIgMChg2pBvmVpxn+KrTT6RsqO84ri+y2t97d/Rj5UY
gid1hb5pUbq3BeivskBrGqwhmbFgGLR5cQinUVImGDYVozFsfmXFEdfSLP+lrQgm/LdNXv3NsG4g
Rnj/gB8j44bxDU+T+EvNYxTL+3HUDZTvyg8UjL03ZrdmJfI/6ZxJnLF7KSKdorFOw2BaOdwEw3B7
oLO8owmEUAecVNYzQjKo5iwrUOfopDPfub7oVHbolYrfTnle2dmv1/j7+M/ssa8EM0zxnF+oNpdZ
5aQVxJkY6FtlDRsUL67LlwX7wp5wY4T8FAnk+QJK8cPEYwfAAMp27a1GYxdQbBv7t5NmpZks6UvL
uZmB/xMywb2Qd2ZK2wIczjSMxzOkyfPtqTXIuLQ1iYpuh1s0uRd6h9O19m1K5Pa9W1A3kAKrIGBn
9yarBz5pq17dvsL2Pff1kcrTxAh5H0O01NXwYY5NuRd4inn8G5M+cBM1j3pzoiYseNxkKMZdR1D0
EUU6GA/m3KAJBX613HgcdkJL6bnw4Uni+qxowVqTtygDjO+NEYafZKz+RbaZehQIPvvDXPnxQwFU
EyJ9TOhBW6ICsmdfJZJYbMuJ4OHaoXTKNC+Jmml53iW2rmEahkJUzfoCe55xa5H6gjb4koVCCDwd
rN6R5virSF/ytzeYZGUs+3E0XBxQJFmxm1p6GKCs/gPxpngUxVqJ7Mzv3ZuArqlSJ0X/kt9vshRU
IqNBqlDMyPcCfpO0Y/4uTeGBzohQe/9QNruY1DBZtPPTfeKhAGSpDKUDgs/I0TWUK2VQ0N2K09xp
sqljD42gD2UZJQSJHXmorVev8XGleSBRn+v8djbnpTlmUpdqXf/GhJLJiCp9BqcJWCvl5I6FX2K3
TC7vLlai0dMX3uJruP7uI8FmuyGYTTxjc7RcuckWPBmCquaQDZWmehuEOQ0HIgbf1NTQ88WQn5FR
ocMI/myrxTCaJYZuqcU7dGJQvzJem9C3qI2ixctNrL1U62CB7caI0A+MH6nQbP+V3+c0fXu/By5c
Bm6DOzKYKqI4TFRgdXEjaT6+CPCLWKps9ZuxIjnKsd1G9cpNsh/VUPxWiAp3rQIjShNDC3UJtBis
xPR7cqu0yTM2g4unnQDEhcpBlSuXvIGjBBra6VBYlYztITzju1vPwDWe/VLrKZZEculNkoSWSCIR
nD/gLw4Zs5z1U/HWoshIFmrhFyYX9AMDK08UmFhrkK2Dmb6pzLH/NwpbHaIgYaYlZycuVxfQeb0Q
vyB287gji7hnT7NKDPMJFWoKZ2TN6tGAvYZVAwDXtd4D19wPx4DucrmzC5gGsI5F4G+FpljT9NoY
77MIc8XlYVHcNYpFiApPjs+jasQEPCMwSWvcQwm0anVUO7VW1igBz4KDql4aQ97TAnXhmHhGuATY
LOeRlHnuTtG2YFw8jMRQquJD8LnmD3bjtekL9xGydxIM2hCKy24AyqFFQr3mgEf76rL+BSrrT7o2
O4uEUZBkfXYFbBusbvtOoqzPGXSVnyvOe3+rdifnZ4hn53Ecipq1IFrBHvqJ9p8RHjOUhTKB0G6Y
S+kAyredZjFAvgTekfHOhRHDyv2U9LRYGyVjmGWa8GOHC4hZZoSAly6Us4h1utfysOvd3FVv3E3V
6hzxvvBgZGkcI/fED5adMy7N7UlMgg6Zl5IgGEg4oU6SQ4E5pqRt37Lktr/FcqtXNeYnftCoiwuI
lrPSNSgm2MnXTo74W5zo9yWhCGuk0idnLox2erMrP7BGj7CV3igTr2/LbY8gZsLeUJcVgcc1z0hI
AClLV2BnLtKes3224hBaxgNW65S4d0MwivX4DEKv8JlSzf59hN6+UbUtEoSO6prvYNZ0XG0NUBue
vSBjRXACRRYEI3+RphV9De4ZyNBMoqwzO8sSoFVebzZ++A26CFa9ZXXxdPhEQwHDzy2xgVtaRJHN
CaaiP2NyNHAjixtmUp+dqpoF70q7iiBzq+J32iURYe1INrYornOru1cuRbBtAl9HIka5Yy9Hu8af
uzlWtDKANWcScu4A1Y3hgtkIjmzWg4VRW/fEBYHO09v1BhH5gyUodAhdNJZJzQKxQMCraYihNeip
KU0axkTD3NNy7WZ1B/ztbddgY1W9ZMv3TI869I65ZTp/femWkPpTgtnxBfuFbijRteS5gC9xFri4
nrCLQ4Zgek3BAZkL81sK8d6hIIzEZgdTerY42VEzParSrdVkzSunlLESoQ86cc5PQnlFK2xa7Cyu
59RWdahThF8duQEoRZNmVxyaJvgpF7ifL/8R+ukDtHpd4aYYTm5BnsmHCf3dNIyAniUNZU5IS3MS
ammUKLciDrR3fqglp+Wg4bhQ5RB6w8CcZCEU9Bc4OlSi9oZR9vphPMzDv07/VEmy34W/j2bFl4eM
aNZ7Wb80PcuLdjo3R10UJ8Kr494RzkjeIEpqlQ4GBOqmz05zo+0Hi/B/w4tBazPorRY/hrlplPly
vSN6M7Hs2XOxPy0+dSr95EmkklMoJXGShP3dbzanhQ39K1ebCV1nP9zb/fTyNvoVbfb2b38BTSH7
ugNRayGnCc+rQ1OEnYeQFFj8JTQNjJVZu0v6tNvxKAgLGlkq2Cts3+dxSpb29TPck7X8d+WwfBOY
fVl1uiavebQ3kTOPWo4D2gLt4eDhdHV2I2QlrRSzNhuGGs3w0rg+toFYFHzWQ9+x/WB0c9NqTpM3
9H7LE5Fgf6bKDHN4e5PWAx+M1utVIC/Nfgk0rkQPfX9o9DhzGL2kfbbh+TbLOhcBzfrV5T7hEwhM
rf9tRqE2XxKeCOxRKRp0Y8P64teEYtlG9bD7/EPdSRZBuiOYpDtOiaYSOzDIoEwHiP+NnH4/+FPh
4fKTI9gHmLddFXHBGPlFUHTJtz7w0QyDRU12XbMjmaZTOEZh78unl+KyWFcUrYsi+325kG1wSref
goJVtwzrM2ML65v5mN/lyrrDZHzEYcewSQKH6MDbPbCSYm8rXCwQhdGyUDR6Vz2LdFH38Isq22Lf
US+Px9i9aH4iF8/zynaiKhBKJDwINNmc3e8ovc78OUdQ9jxxTO+j2vYYA0Z95LqMGEoc9JjcFP1Q
n8KtnLEFn9tWxHOMTR1Jcg05p5lHXMglAPcNAgByMvTq+uutCWaIXy/qWNXLSpkpsWwhUnLcYNUp
PCVgAqIomLSmDsSKh0dvsy2Z6VEUTFClF+QYDuGD6DdCZwCLfAV78Rl+gvCA1wzXjtRIzJ217VcB
r65gp9H+XIcJB7t6mXg4LkYiusosLvzmltP4UStT5JxGZQXbBeA9PeDTJrlzXtB3sqj9lExA8DrY
SUIY8O5edmno/A8u1K4IDfeZ12dnPvsEBbQQFd5uX5TepybT1wevzCYJM0KvmZcHGAnwy2fLqbFg
oR+bVqTRp94Q54wiWJhZSYnyqTb5rBKuDAFuYHyvddnkibmPlIzIgOxPQeEYEO5sOldEhQ/1Pm86
CHgCLJEGpC7vQelJwSa11KaG70XH7qYmdebPcXM6xCpTpQOfWq7pSNU2FnVQvj+InT30jFNxRyLk
JuKPDFum2mf07wrfMVEk1OcT8RisZCPTuGskAT/VqS0rr9xIobKVtcIPkViCdy6xLc5pnN3udCKB
9Gjfrh4epxf9ilJcal7cT8U6SD4DeMVLl4Z/iqXlBRJ8P/+PRW3x3kkUXdAqfZodJuiwYkVW3cXg
7YlfXuUDKzVV4OHVlzJzoSlvSlmF1n9yGyF9nKSWxFDFXxgaCRjRHkIfGs5ThojLeTf5Oa20DqCb
WbVgqPdWhZAIWqQ33IOilKirjwSDfmPfx/MSgNT9ISN2Qbi956mWymWKHXordn3k+ktBKlyn1iGT
xxgGsYeMFonNV3RO/BAWotgYJk6n4wp1T/+5Cb27tIc2ct//48uuNQqRRiBYxOG0JQsbmoC7m0Pe
ieWW8gsNyBGwNYXVoeSyogChULjkLXnoEiSyNMgBoUoEGHWqWbv8nvEK8ZEWHPtFauXjLA2ju3ZV
gWGf5m49olurseWPZoq5pRpERkvqH+9ai/XkQI5mx6lSiHWICq7E/ltTSvV4LuMWTA5KGu/8cfoV
f/i6iJkmFg+RlsFHzCnjUwhiM9txsk/OTj2zpAFMF71WpzY7Qhjz1AnyRGAxkRATTTNizTP/brd1
XFhTWjxnjfHCiFScaNhPnCKvVAG5oPqpVBAhj5s8f8SppI6oAAkySfy1vaAFpC9jTFh3vlfhpV0j
Me2w4I0Dxb1wiGSDE0amDvigcVkGQw4edNAZPgoAIwPl57+NB6XRS3Yj1YNzH7e5aP7SAwvGPfhj
o3e0htJvVoJ9YzULL3T1oeqKpHdJDmVX1fAO/5No8q2HzRPJUKqA1O4vTKJ6NrSflRy8DVFfAgFY
e98pPlJ1DVofxgp+ggc2Pax/3lBqGK1XmupiYKQYuD5Ka2TqSrrrdFr7enJcbsymcQog9Hm6kpsk
Ysg6HAyJA6j5oPdPmAkAz5EJOL1dqXUpTFQY4Zk9pPtIEIPgsd1pBFGAMOjqFDCgjWRK5tTYuU90
bCcQ5cboABeBuYSF0VKHwWWdaDJY7iZUktAx/JXGr4rdFyeQrVISM6et2Mtnz/ilfGaZmhzglP/Y
MK7cOdFeZI7eHfprFBmVmMxkF/j0bG0YNB66QIFjBXMw/yfoZ6+4vIfWhWEl/C0uBgySkKIFCDsh
qfa/MNnPkQVOzkb4wH1Yo8AZSWQ2Q5fRXbLP6BEW02ZtFr7wPfl0drnX67uvf/4TBJYyEY8ZNjYj
VP+mjLVwkO+irEiT8GrEpyfpg0h543xuFJDwuBSAU8SrwZbpZ2AhhfILo+6TcugG8qGTyCQ68wDR
ZdS/1tS6/ZleqhtOW2aJ2Il0nGtgOIecjQEa3dOl5fu+2p5Jh3RPZahotyb25k6lEKTUuilaXJl5
OHMqQ1AimXu57oKXY8aIChla8a5jbgf34+SOnllLRx2bCdmI2SAxN+Jx4A4iRSjvMfB2lNTcA6v5
b+RebaIS9SLizCVQFIJw0d/K4DxJOqj1DmDUYmL/0xphf8TOfclyLF+AgRlZ3uyekrxSfLFguKwz
5Bb4LGW+YEmnydVdJLOgtBTZzqPl321ITT4AiH8RJHr063giKPH6D6NcmRdYrP1HFFRE9Ri5KTzr
RLdBLpcTxksxyA9hQOxERx6mQNI90uEx2FtX4+L3DUKN+FDC32FGJPAuke2KCchl5hHbo+SibdMa
BApG35V/0g7IhRTTTC9N6uQ8+L7ybk5lLoa6zLT0ZjtjVMJwvSfmY6mekWA7hhcApBs3aIRy1bUm
LsY5REAfJX84iPbd6nSdt0YtDtMNIb3oV1ngcj1GgT8xWo0NJeIaFwX4hXb22Y5J728U60BJ6rDd
Wu/mQULj0aA9xpYYIhZLeGGlGTQrgm/DY9rcVRJgihKFyNbs4EyLint7b7doiS/bkJKGBx1wquUw
eHwPFuTn3hho+yqcQjEPPQDdiTI1ZGFiX2Sn3a/YBTmgCqLZzvc1OWFgU6ISlfdC7MTKEEeBPdsD
/OmdQf1ajXkHBj1VTKR4qRNzmftJSS2c9/h42yZvj/OJxAvEdb3fyPdhkCVy22kYkmuLY8T8/2VA
Mt5yJ/pFGtUTVH5f3rTx9QHJsZ6waWXzJOJt5hjvwFfy8Jgz0mQUKRdSV4zJAsMbqh1g5sEHvKw8
IyhkykUWoUOKj0hSC+Ydxy6CkWr8LnvAKi04w0n3jNZ8PqtIjICujkV9cj8neqBVSUfr3SMJ0Y7r
lvSedfHJiQWONZ/zs+4dtDPu2rndeDtwZbRa2VAu/K7+fzBGTsihabClynZB+UnHlkJQkF6sriMI
WHixCzgquPWPQzUYKILNfQpO96yvLnWbQvbjqDdEAVrBOuJQ1B36sIkwsEwq9m3I3L6fodAstwzm
ue7LvtB9uLuDGR8sBINcs8OodSn1UnKgg6xquf4c0nu0XvGTHrc374mtq+LgwvReMhhBIBKVNM3m
8t8lrHa6vrOxEzF4k0rJDEyBELDafDVKgWs7NG5nxkyxaCbJkOFAubh+u4jtB63d+DeBUfhVww3y
76bsiVtZkLzGJ6cExY5OY/+4/LeSlR0EZMtlO7Y7IPP7uAJFrkh8UcPHgag2Df1OeYliugDXLJfu
msjkz+NBdjJG481bh6nDPGsKzmjmqexys1AzEx7+exUp+U7RcHIeMk/BEsXcOA6kRCb+GPvfI4Kh
KBm95eFDSqd6JxVjX+Q3iN0sX4Y/Hpw80Rn9IyzhFpXpZcI/A1/28iLDP9hVuyljS9aMMDHthZiN
DyY+O5eYpl0UBizxp43Gc0e/Lj7iezhZA6IpsMyIx0GMBP4C0ab+6R2khXVTd5+mCsI1Zub9LRV8
3PmV/lQM02/o4FSI8x8EOf7SDy6sRlh6gP5On0flyRpNGA6ZCqmlmu4Ds+SGaPhm9d/FC9iBplj/
hB4PfafDoPAufwT8cpeIZ/v/Ku4OrOhjw0BVpP0aLfYpmnn/CJZ0WG6A+/o2E94ve2C+5t4neqXV
YbvW9L2HHdyESsY3FG++usAgCteoIPRsGOAJ8Km2tUFtdjJhdPz4Bp5Pzyz+9erjX0j50NDodFQI
VlOa0DNyub1CEXTEFMTNWfJwpDk7N4pNZ4efHXdswQGEEepraLNpe6sun4E0ETpCqBDC1vhEliyK
YJwLC31wMKBKrf2OEzn+la0+nXI8V5o+71pyn+IDiuCGdE+6fq5HhW5vPHM26uoXSD3MU0sqLBAl
vJK7ui8c1uNPrtU4lK6AjKit0AOxPU24QK8XzOd00IfuDmr9EXamKYgbMq+3IglyLDT0pZ/ufZoz
ZU12RlbO32DJRgItR/HvBC9PzRQFW18VxfLzBIKI8Hv1S3WF4L8pQ54hTFd0YFeL1Nkvtb8qgWY2
cBVohGtP/lXOwzwIZOpJWnTINCtjZGt4w4sYnuGJ72GKB2yN7jqjAJmpWtqFGNCnjcwHFf3i1xji
5bO/wuVueMT1xsrk1HiMv4TPAjNv3KscvuwGQAOXD0LBm6sICjNw3mlEwAAHyVXauk3ipdoz1Lv9
IyiayhxtEPgd2z9oG6Yef/E9ULVc+80NLTl3g0DewXfitIBKzNNseZHj0WRpz1DpfEXWJhvjao9I
rdGltKaBn+6VrXUBJhFNltqmkxsa+jA98cHD5ErpabP2FmcdQKbWcvnsuTV4boYZLi7K2tINhESB
P2MzcqDiN1uvpFVVSDYQZFJTMOb2DMYZNfKPW0Wgr9Qls4QBKz963JS8nwHgvWvjLIOu+UaoVCi/
Nsuyvf2KG9IdOIXpjXTKVH5NLPAmD4TQ3PJ4eBkCbEtJJ7oAyRhT3E456+44OJGNFi+QjQIlMix8
S0ANlg5FLPBWkDwEBar/iUVqiPz8Hj71pgoEGhLim7bNt4IKzQba/fOPn3bc94LCw6p6w2TJYqi2
5DGXrjBD2QllPkhvyyU+u6uJSh1PgSM8yjstTB40ovJAkfQ58/MnkIDBhD/sZ+TosPnGzXGPoEmG
zAtx+tljVM77cQmfiMViubP4Nqyr0PHL/JsAmpCDtdIM+xYaQJt/+9qoEuhp/H6DlSjz2QjQJD/5
UF8JaAY5DUU/DSDd3gill1U6u5Wjz298o/jzKgj1x2LcP/CDLWvagLcmljExKcohWZ7YaDhUEYZA
4Gsf/mrA38cdzXhEPMQGcaTKJe7IJap0pmvrnDT08ZcXYxQUd/NqI1bOKWbV4f7nY5Qfz3HKxVhb
imvhcJtXudi57V6LAqBBVhccIejgO7RvpoysB6mCa62rUGtlZLgWQpkkVdEkKh9OxZskeW3eiIcj
6amAep5spX75GByo+gvPFYmT5C4kMqVQdGPM8/eBVrE8+xUlt32Rz3+7NwTL3H66HJthC0B2lL6+
7pOwRF2zz96IvbLnq3UiMYkY0v9TCONnYOUd/toydF02aI3+Xx/NTl+8vLlo1QjUWIHRm0DP8bPQ
mnTXIcfhwuOwHFK5cs5I51YD3HIYitRXcHr26f/6KMyxpCLedkiHsgw1nxzoHBiiQ0zqzlbHJiKH
iJBtGtQUGs9hw5CpHcfntKXgZscJl5zGz7VA7R6jkXJkxkGn4xwoPew13xDso3r35o+tXBkd1wsy
OlsD8L/v4FIFlQT9MzPiD2/1w+Rup5Ae8hzVR2aY8mByDsz4K7o9RH2FiCW7ozPDE7bFNetPco1I
0TINiu4dS6hfNipaXj89Xls9AXh71jfK8lvOXtZOAySlzInMiVCGMqE3V7Q+Vhbu4j932DhOisTH
3Yt3AUiL50zi7bAR9i5h8GbiqdMVJIW2MqjJLV84UgElRXlGgglBz9UqRW/NMWvfNxaLXqaD3qhn
KUmNjCzpxDxm4C9nHMwJ/kJ7fpKtCcCv8N3/GBNOenO2S4Vel+Fjxrx4zGg7hYbvPFug10f4Nchr
cBMpTtxyVmeT/aOVISCr4FWTHpsebRZrLYrZNGxmv7gOM19vGtnOVQ0PrJTCow+vRJCakYtEhW9K
bMNs0itde5cFftFRWuUjwEV2WMf6S5NpIlwrSjaexwB7xNuGXUWfMYcDo4ZMX2PWiYGgHjYzngza
3L5b/Qp3mRC7iF91KoTnkFqJV+L9hNzcE1b0Eqx8omDdHuUZAYe0Gsgp6NihzGyNxzFzdsO5H0vq
DZAxbV2idxOyChQXIhEQJ1tHq+7thVAt3OGH+7lYOqzeVpEHMCiGdc3YkZ2nEuYFyXp9VfCM5YYK
TzW//h7BkRuzsXZeNBoU9YATZolmdqjknLnJ4o1kwtQb0UaRVxR2J0eVrEDiu1g6+7qnHhP4tkhD
jxG1Rza9ob6MCuMzsFNWqWLOXmIt1ORtTKKpTbBBJ4C9bgbPrx60/Yq9R+Gxgm70q/2EkBOxRr0d
3vI3E9yXbJVrfdyGKjJH9QQDv4Kf1j5284iV8s2FpibLiTpx15Ud1mOR6rRvNxXBy6ZpTe9XLj2r
a6SWa6DWtPRBzOg0v76RZqz3XYrPo1MVNmhb9e616Jr1V/88tes9gANz8/NkSf9LLBiXkbOQbHCe
DH+aK/5AEfFS597vxLJvcyXZgpPUfkUP0v6oIwauDKxpWdcgT85IPtAiLh/6lDe94DT4bTAt/5wo
zkQWvG1X6rvDGIVajYQE6Qs64LEbgQRubPPOd290TS7G5W0EOi4BQnt2Z+68lYXGV15asDlHuMne
qzuO2jPqa9UFAAD0GN825tn2kvDcTTm7BiT0R+xFAj4+qrNXriERRHu/AaM+5kgkjzHmGPXx+QN1
N9aEnqUBj17E4IHJZdegoQLRBemVjofvdWU731nnVe0lr6e6zIBBfiWetdVds3DpBG2tW/7mX56i
xGTw/0jJOAXh5YH8vMubA/DUog4GQS71rQ8hEa6Bw8dHEvh9xZsUK2xxEe1nx7ftxSEjzINdQrbk
4PAMmd4NO75siLtZoky/eYb8L5Wny0fSTuvcDEUg3Thp7BlHBPqmASxtEMrZvBs0X3k9wRrkLgXC
RrxwMKHLND8oiQNq51xlo4BbxuNer0pzwxW9vXCvsGeHXg4AyfnSiPiD17WMXhCdnCrC/PJBPcn8
M3ajjEWjAogSRxAWPfcTmXE/5NcY3H3HBFRoeeXzyeo9splii0BY4AIIQuaYCwcSm0/boA2qRGP7
MFI9GfU5maJ6y7Fgla5FsNj61Oo+TdPq657+W/SVRAUnr1SR9JIHe+wBnPl7DZu3xvnzUJafxfym
LPWNsZ/GSa2SDs7Wc7/4PvV/+8QKR8iY//VKPNQ33acq4NMK0YdZCbAb9r83R2v3Rrxs6F8LgKS+
foyBcrHarkVq199fRgJKUG+mMLzsChANdmKGLIHbTS/vzyDbs17pQZ4mzotBdXVs2dHHr9aLl9Yb
1ASjSpEv29mb78YK7YXyQ8crqpaAyVq2zwxurEbdHVGU2j8nXmY+yOjKA347DFO+Ak37hcogLC7m
P1COYH6Zw6xNjdW/QCJy+NUJMjflTqo1Lah5m7bVfQSb1OmXh3hpAgjH2KrSauYKBR25DOZK+qIP
+ykqe3kWcdxlUeQYNBSlQ+axU/moFlEk5vPOqcU60nNWJ0nP4P6uLKbfLc5zLgTdvTtC9VvhxKg5
FdRiOSX0DiFaIRZBJnHMv2eC4sKZ7AH2pzB34Ouxh67g57oas8s/G+H/2PC9FjHlG9rvb2y/vKji
ldUTyoFpCLSV5gGu3NfRM1PMb4ByuBS3dd8eayWSJqQ81r4ZFLwm0DwKSGUjgQze8Z3op+qoANbi
rJkFgoExSF/6vRBOCt+d8Shh5VJM6Ku+sHOTQIaGwoPGh7HUgtJ9j6ZepX3ZASTzenE/vOV3YWjQ
Apl1UiCNkqedBB4u5qCmQ8TQEOb+W+9x2fWYWj8OO54bd+bNTu8MvaBIv8eyp6GokNc6QJiyjvIo
Y3uPfxqWdfgeLMaY52Nd0gwiqunwKQeYfloWpfBhYdsuUSqUDnMPhG0u9vVR/TIhlhwPNUpe7Us8
FNzXP/ytpadBcaZxHNQ1+rZbEdSo3jVmrDa5jtUOlWKe1UNCzRO1cm7Fzl72XAix/ts1h/ayy4oU
fVjFe7mi9IzloDQd3s6AfLMpKwwBQPVWRQ+27Xc0C9xpjU/tWZgZ+N+jKJq1IsSaixvImmS3k97R
EjHgY1M3qcb04XWaImzwoIl8cdUmTG/m76yP4ZXPPyH/dmWuvjPP5N0iLrcyPGvA2NDTfddMggEf
O6de/l8SgFQukageEuG3PWLGTIyzlyTrHHlUp0XKzaZu/bbm9kbiz+zGY6rX9nU54ITfBYKzfHT0
IoFlQLyGoLQ07vJAkK6FjkRvIRFdIZgxg126z7Ctupm9k04+Ex9THAx4al5fTJJKCFrjPFLuNvSN
3MjaxUAcrlpV1lgEcNz2bklvQn6jP5pDkL9YUzkVGiFpiE3h9EnPXQAR8w6+yHXU3lAO1czx6jZ/
bEbv5r+isDw3toEzw8OIUOYe/XQPtUHD+7COqtUXlN7ywZqviXqcYCXB7+YFHplf7lEpyqla9+e+
ER+7BIYNlH1+wx9TzGeJelg+GcidlhIj9+pVy+VL9ej13YMAnCsuZcv5jUM43NHRPN792dcK8h1M
SK25/i6QPw3Ey2uin1r/iPgk6itZ9l4DRzeLFyc5VsV//6p8gHjAl/hrrifZWj5v6uK9j/Erf0tx
ujl4geSOy16uiKxRu7yCdy4HDgCMSEHsjyg5LSrhyq+bRTjS47w/TjzO1Kf2ud8usZ6i7zZXMYPM
9yATn46Ai++wAOrYVW+skfO6PbyImdqaAEV8xY4OcXuOddpZNbsZ0tK99RAjNUJqzkHfmcxM8B/y
HUt5gs2NDmz99vgJl6VcNp1Ubo3IC32XiozLdYW3psOqYRae1M6ni5y/7yGKJau3LhMCwv117Ca2
YZSP3JKQKfdhTTfdafj3eRQNQ/UIwgJO4hMo6v+J6JA1l/NnRHBaGJ91UcIP2Zt+3deno6xcVgWW
fk2gS7NgZ0Eg+GEePbQc0EESuYY90ifrxowedikKxosqK0qJ21QSX7Hb/DSE58XeQ2a8gNRSNrAX
dLm0BzypkafTliYgliKRMrrZhjPa4ON5s0dR3QytBUmo4f+3L3FYGNs0yip0Bz4IzkC+l98h1Ii4
DIWTtqYMg7bGvBMHR6tnU2V3+QqmNs/b1M3s0yJ00RxvKajIMz+tt3Ruexm57MLE12ZZj1NqEFKO
lpAdjp9jyDNDpqexnRBxh4SZ6mFxgodaUAMfaN4oY6zi2pvh3ZzurGQNsaTk7f6Tw6g/nnTCGWl0
rjjhYVJ1Xl2xk9XPJ0iDjK32Qj0ZLQgSPYDzC+o302DJWccTWdmvwA8ETDQxvEqV0iL9xG4V5Ftb
04zZQVdVeOvzBuKOIDCC5+yRV7CXD7SLadp0awB6Ja00/WDq1FFLteU70udlbqro8O7UEuAqsa24
P/fHP0Oa/fDviEv4vqNfVuLSXfkhu/hvvYFi12Jx6ozW3rjjGApYfbkZTrcfC4xS4v3B6XwNJ/V0
iJkx2qPUmv9vYRpwbYr+YZ6WJ6OfVMQUI2nebduWdWWMqAIX0+d59vsxGk/a2FeSkQM/Xv8HaH5V
vwHrpBzcI3UNh+7MRG5zZhhDkoQJ8f+SE0/H+VTSXP3hdQF80Q6IXTUEctXO9Xn73OPgMhEBhPzY
5Po4ebzeSFwUG3KtwHv9AcduGTajS3aXafmHu+QEJKeJ5GA+LEXJBuSTodXnvSR1SUnb/4kLh8Gp
auqQcDRNu7qoUiaQwD0rVPsa2bHXm88pQJqs4vAZDx5bMf+DSXt0hyqy9i4l7JuVtXja6ikVbbcN
ZKNxF1M7XZAmCoJal5+4O3KJcegugB8LWvQQohdnuUXfSAlVA6451krP3fUFa9upM7RxM/3DUN5p
Cw6/c/+NPU7nSx4gjWTf8/M6MXmwmvzhQFC43ijL8kzWYCzprA0v3HB87fDvBpVfhRPZC9RjQbGc
0py9fv5fetN6RUyomKhm6/Mv2znCszxTKIVLFBAFPs4F0daUAuH55S5lTHFUE9N4WR/tRZ6ZfekT
eIQ7mXBcuXIZJLqfxzwkDSNGY+IisNl2/r1nnWsMQcYLcgOykhpi75y5SQ6Bz2GiIukNFFFfb7Ru
J1g6AhIsrC/zIc4XFJ1/aC3+IbYLs577cihGtRQdyPybBJtk8OiS+1Ze1UuG6D84B8Pg4/F9La21
OGInjJoYqDfgwPJ5Z0e1UabYLsHm2PKFEMN4UUKLOAKj+sTY7PehVvUCJOTSe5mGsm9ZkH7J9+kd
UfRUISko5Q+AexfgFiRQy2f+GJZcF6trNiMFoP9cGb6gajYCIF64++8DLnWFRrd0YXjD6VFLkfXt
T14XNh2JNk38yDXrZ0nznI6i0ZZwvglfnuP7Azar7O3KNN+vlHUu26ggMkXWLLn1Yr950A9vPlZb
wvnGfk6c4wUmMzf7AgIQddNGDEzzCl8NjsiJPc1yp8tGVxYwO5/fiBLi38/13lXBgRg48rGyMr+8
kDj8xbPuPZ2WTL5zJtG+5tG6QVWtxabz4yTMAaEyMHpUwTn6mL9sKYzhHi0BdhAnWWPMiD/Mut1p
Q/DHcWx8ZHi4n4bSmcgUKSXqMMHi+0Q6Rx7t/6mROW0Wgwa4mbx5c1m8Q/xXZF7TbCizEowLBxaL
lhIdtczxIUUWxZcRjcdDnoeMFwCMRHEsRgUwmXPn5iuqAyUhYlT4Cm/XTkdbvM07Pc6rBHkPLPIi
J1fO6Zi3yKDvwzjG2aKMALEA4wbN1VFHbxi/ItpIR49ezJJAha/MIVnn1zSs7K0e+FnchDuwlu8n
DJd8q9RwxlqUCpqkPmrcYve0J52OB/DCMoyCa7C64tS17UZetl6f4N5Ipk9iSCIA1mdAkDjc10JM
bHNziohx3KkTU5FX7HSpCBuhVpoGJwS5pbSS7KF89xq7fVpz2ynrwMjrg/m0QyORE81yaSXGhQpl
p3H8fomDK2tR6N+XUHtqsrCHxQLfPRF8ZAl0/pLDYnqrfuKZpUOAmvT77n3VuzrAlJX40lC65XZf
6PBh3OBNLhWuNP3MgXyLdoq+vM3CI2FguhLjhIfKsfyZJ13wZWW8b7XpZTR2282SjP+Mf84RoDsa
3ZeU7QyPPu+r8alSadvFdexM7LpxwmLoTm3iFP8ZIpRdI9lB3Z4xiYXJGAgriAb9loUN3BwoYrLa
KStk6S5BPdtjX4ZtIJ2mAei3CoqW8+8iyxvATAozqNiPc6c2TqQyYtxw4GJgsbqMkm/0CYQQShMU
2bDQe0aKvgSWS5Oo9K4AM/IimWtzfkO+DskbqKIy2LOWit4igP7VWxAmuvPBFglmR1TGA946g4cg
v65TV4UjND7JEe0J7I1qX6SmrF6aomrubJw4EWiVUg3zSBUddYNNu0BsVhKV+xj21QVMfJtVFP+S
CQj34fIU+nVlLXiJeJrFpsw9S2cxLMxWhlvu6GU7dG2vy9pJ2lYfbf/JG6ATFCCplEc1z7Jv9lC7
XFYQA79h+8L9mxGuKHPE5X5ogrgUYlm/5UmUOmj7uXqEmrsMm7mA0pKiumT0Rz3fdJgeQ/u4hxqx
25b5ZYxHohxLWrZCAXu8H0Et0nc2okDENPZSrfJ02vj3dJsNdzU/odLYdjxd+HOCA+Ys/RmfNcu1
iUfTcUMd/gIX0ubZUubOY/zornSa8w9ANU77shybuU25pwVEVW98ui4i0mqEOASvKPZ7tgMFMnIl
l9wwwuz9E4EWyBPHXJYZCVucIEHtOAkIJjqGMQdzuv5Cm7Ps3/Laba88Z+Hn7t4nVZ2C15TmLNeL
BwcWpTChpUvo+OY0iWtxgPjXefqFWFTqtbYtidRuQnYil7v9SdDlPx195aVB1WR/WARzZzwuqtg+
nCY4zbPvDbbjx3aoUTPO5BMBMxzZJcxnSDUmukGga+tM1pspb+1RRkQnPDa0PAkj/+oFRjMLvjVc
RXOoFxCYs6UAIOg/hTvAR6G9TpjVIJiDeAw7qB0Q9BL65M4bi4L7XfPWfIBPwdvrwe3r/+jc5lUM
nyt4o2y5mg7TjOI5TQshc+magUHnOBgoT5QyAAfhgbfzkgu+5+dgFSa+eOwq2dSEt6PODUMhlZDH
QeUJW+2gL9QGPiFkHn3arkNrSl8xHCfuglANjBk+V1FQ/Am43Me64hWVhoiy7r2GO/7uZzXjS4H2
yDhdCJnhC0zDnPWN0XR+fLoCzGbpIzRijRMkTBzaphnJH9snFFw7sChyB1vMQFxHKA5UNmhsQs/8
11KQcdQd6AIuu3jaUXSz3bpfdwsl0pT/3JDKlOc5Gm/jiFKwLhW4VLjM8ovrypF6AkN/M5ynt0W+
rhP3sqz/xQFbdMqrEpByHFpL2guZn/D0WmXcnVgPlOP1RSTA7DxGLIHeVso+ykPTRj+vWJqPEmzd
XZja2gvKUbI8nQcmO0cNrgbF6v0bp9O06RpIOVecwcrftKiLS5O0k7QjnlJWf0daP2r1cv/3NZNW
rH0JYADmSXWGCzN5ej0sPiSfRNxgaxc5iixvc+3lnuwvwSiRmwKJuZuxGifWQ1bfeiZWHoMGb3ov
zZ37j3EFTGtA8ZKZDVKtpLkU+vbdfGDggRJRmg/LK0mEFrf+NGb8/rqhj3Xd7y3txuddf88Vf9+B
jQtCK98uJc4y0Z8Rv2bxSxLayetDQrNK3v6fO6RrvtZtSE39GtaAjPfStAbMGW+tG3ECEQqbyWp9
vkCwzEusKSItwSDmwlJ/HLyPAJ4vmfcAW7GflGXIz0WMbu/oRTD0O7dxyoVHlYRiWPNeO0KooWC5
4t0POPqKPQCt6wb0cdbIAwbUaJ22Fxs+ZEoLKXx4rfiHC1jhM9PKoGZe3zD9FZ5yD5nBy9nFP8u7
MbtFGGMlDqaoJQ7WMTTixhrN+ifie9EeUUpqXB/wicVpJKx+RMbvJrwflc/o1cDWdZDDpFnypeQx
9WQ9BQXSslzPuX7xa+FO0wtZ25gvGfVD/6tVWCFXjUmFpTIBB68+YCiLxepolnfQ1xlLTRaspc56
W6S3P/MdF0tI1+yB6XkDvVWTepG5w+C144X5AYZZyhzWE6zJP6VvBxrhJfzitFUUqKRQ/1oJwG/Y
nFhT8QVav5S//CmDKTRX7uSv5viAeICB6QlPKnNTKqsX+eQa51KBhCM/1eYesG9NeetZOZm57Dzq
K1gL9TIsK+TszbxhnmdZ9ybLPuWZwcd0mYVomn7SumzJgyoQrSzIIaQovSopiz8dg2N7qDzfkBRt
zyeJhqq4hQH+QyssyUJ11pUBGG8TlZMfje4QufVlSJU2Fs4Bo1TKt1gLJj1WjWVA9cI7ibXBVvXs
nMMSNToAHyO9qrOMbLcSgWVSOZBm0xaIo4J3IgZdsPDKV0zfTmgy9TTcLhiLEOr0woiAT1DwVfCq
kGzNgx1wtsdjwxxZQd78fRxgEHvhSJN69pJ8iwRO/D3CrI35rDdpxODwgfWzCtD0Mv+VbJFBwcJn
xNbskRi4EyEAF0/NMmheEuJri6B6rvetkxLQSpXUcPhDE+pRfIINP3lmPtz06D3gDfvZu2fc5IjE
LgY/MX2KgnKXbe/BXIn9w+1kT1Mso5uLcFREGoj+9vKFBuj4TWjastPBO8+EjMLTBE9R9E7CttIz
W7Zs64TdpqqTdcaOPL0QANfjLXwCJZz37sYJiBDHRv0orYMlsH869iS0V69NdT2fomZLFBybobmy
sGvpZtJyE1/PEfbpbFxVkeZEQrn5meulwa3q3hSX5xi66NMTEUxKVzVkwpCfsv52Oc4P1HcVccpF
dLDISLA2iUf1StH3gGFixtPSjqNvAfujbuja0RzPvSiChzLaYfjQpPWQ4YJtMtxKC8cXLJqFMI73
JDF1u/SrBbsnviI9h/zpyx81qqmGtrop9akUna8z6Djtk9di26NwO9+dXY4ieqUXW3on6/r1jBQp
lmsdnvHtFgqz0vV0M49mx38vFBNMj++eUgaNrJerklD292FxJD+QitbkPayaK207NvqXWSyZNwio
N7+0QJzSCGTzSzKUBr9c9N1EBG0HJJ4QUA+HJzj5jx+eYLwsg5VZESONOnSNjrOy8qR5ShjuV5V5
TnkEHhp0aOYzqJztU9KFJX7HVpDYWjM1BRqBYjVdVuYoi2c1qVQLGCkiNJoofRd0+Ctf9s/eWS1F
fxbquEQq/O/KkFJrf5aP0g1IMpp8Y0vdIFGa8LO1rR912BwfAqTg9AgTLeuh9HNQjKk6ERHW5tRD
s/ty5GroEPHoJkCFslQrsjFn7vowxXt1i/FJ1ICJ1UjTvNBmJQKo828kX7ABK6V0szpnEu/RnZpk
KcmJEyTCIlXfPOWCfWWvqMnMqDFa6ppGqaENa4R9it2y3/LpEZy4sNskEAtsAbwQ34HfA0whrRW6
UzqK0fENXWD5w+K8nrHGPh643Mr1qe1xIF4laIkbLtgKVLv9jmI1UhpaOk4NkidCMnfkQ4JSsRqs
OXT4pvRl7lysbsNM+EUnuAYQZlSI+n8RN1m/UbgxCpv1DgWwjCINpPJHlhaDkqNC68IRfDoRR3QL
861uNdrdT0ucmOKY9HcB1kxYtG8xr8tu7r19ErGzURT+zN8V97HKUHEZn9M0lOGx2sx6JhAACvVO
dCAYWYvE1mjTWvgKDNhfuDuV8CXazLniWKhHQjYeTew2hk5/w1KK5APmB+l/LQUfa7gjr8boTpUv
n08u12o3FfcJTrsMs8Ujvah1KvCVhaK6KdGf3+qM35e9XKfTgtQ4Dq1MG9DGhvJorsB8RneoH3I/
F3Lg2fWGA3m9VaHAiJzhgIc2i5G5nfu1Uc1aBIuQZjGmK3u6dr6ziq06XZPjB1lsTQwsmTzRRP2/
xLvzTSLqegWkmLKcr/uX9kwxj5pdfHScp2k5GBHcJlVMrwUSQ08Wg+eVbEGtN+bCKDj/5tGwBxEg
nzax4kOhz7pGFlzksWpWQ1JSuvM3nI3JdiswQ6d1k5zhF9ew1lPvdyqrKN3yK4vKDaddA2tu+jC3
chWjjwyihxXVjQpowXWILAYAotimXXS3lmNybzKRlr4f7L/TLBBvMvVWrXM/Od1I8Xg+gbz4D9my
PzXDdCTwMEcWemeN5Wl6dyXBjNjqew5s9gClbE97+ufeN8m+196aozh0NkxKK9i3T4ejp49S3DZ/
Z8y++1RX+JmmHDbR4mzQex1NSZB364LHBn26EFY9IEB0qv7LuluxR6fI3fpMh2GX29TZ+ZsjQLTU
O6YJbKCDJmOyWgQ8MTbYIM9uPt36GCFCO8+tE2fdeJOjn7CMct+v/q2vwOx+z/rRjhSUtrTLjBwo
Qv16zwU1Wy9mzbmSWn9BU7VJ0+Gzk+e7ZIfpYNVF0oXgQ3lErLNYKxlMrTt51oVU26mEsMbtJ7ki
gufg9gz/IwdWhchpk71cXktJkIO3sbZ1sXUF+RBGrpxXutrXigu3rkE/nwBcNKRl/R9dama7u2lk
PJNIdMmOBh54+WD9aesTvx3uYmO1LCCx4Wk6glDqb0ehq4JYLvObSR0XWkqBSBpe87skICGJrtkI
JrGUbwGEUJAHvTuBvkFFpBwMm2gWggSc0b2jl3F6aB/HtGSPcq/5nqtV6R2DUYrbYp4LMdkp0pvc
H4oiKvVzfHaWJQaUnOrptymjCKGMtCQGDv6e6q5pNfQUMUdn38O8L2dD1X/zmRn+Ulnt0NyFcvhE
BhBIxMj5SRDaQOjNQpOXo330jWJX7zz4WOwBDyz6MjEhg1wnm9n9XHo1JvXHC28AnbqtCznXQ3eS
rLexaIdqeXIecJxeMBoQLmLXVxBOR9DWV3tZagdzXXe6NSDbJC1ttV3WHtiLkBoRieLbddFwrbp0
cXBO3mWMpMrvPPAcqAYjjQE4WaoNQ0EfEzSjMWUgXA3e6sGisMYDDHcUQQVlA+OFfyaNNVTVUyl0
DShVl0Tnl+6XoJ8V76JZNbTa8Cv3FYwpqQRB10O+2qH8tnRw2j9vD0CUJDrsWUMD379ypPUvsnUv
FZGaA+NX6LTE+ub05otX2DmSLaX1l7BF6quIeL4PCwxxq5kzsRBB6J0Bipm5dFc2zUOAhJtodMOM
Ia2pTMvMRailRSrn5IQnqgPT08F0j9y8axRjDCXCcchoGL2yUa+GoX73KZxkI3sRy4RPwtUExGVo
GprwvvOQCGNmhmfmNSsjAwqnHaDGnj3yxYUniwRU6FrOn7Nl8TtJfjEdOANehHYL1FLYXsesjQBk
IYrbZxw5sKTCR2otw54w7yy7If4c7kyWHUtPKbz8rlBT6SZMtRRfoQ7kBJ+8Wy8FHvt6Fh2JHOt7
MCuyJ4MjmMEknQhm7GXmeDQBVnSpyF3o9M5j8Q+RR94TXK1H2Lp5x8stDGckb8l4iqHIIyeU8LdN
HuE/twpaCnQWm/O0/jZGjyq/QId0HL3G7FHgwmT+zWNIL5gblcgk7Xzif/PWsMX63un3bckbQ84t
FwtJfJLzSoiSa0mHFeoPXCkkODBQX0JNJ0i4RdJtGHij/LN6Jh/TQtkwsTnupxypE0+2sm2sSSIT
N1a85MgfhOa7yAshwPCIG3Ia/0C7mT6JvZXV1M9b9wSBia1hR8oNv+l1WeAYuCG+6s9Cdx02oPGy
XFNBA/LzHu8YVl0N5MGQKKFrW2SsMBkQORb2FTirFqSI9GPwkrKujZAuZn8SYiXFcIO+dPZW02L/
qraKH0lOqfJR3xU/fGlShLKmfx9IBTSAPkUm+LUuCIvterArdAzcKNDE5UH68EweE/W28TsxSWcG
phR6w0h/oC9txBsoiRyHz+bt+ow3ehjm4jVNkA3OzbKM8rZPR1uWX2fzJu37Q+/WL5PshfA9544c
fk/Wy4KqG+HKfcxWPop5S0AMG/6PFRp3WkQeV9I6m5dWn+CQ3yaz4K4vL90IKuF/sTpS5Yu2wJNU
L8QJgEbJNHoIx03adInZEyAaNaEEPhxyCHazDnnVhMeIc4SYPvFDhSI7zib6aIOPwxjZax12y3tL
b23BMadRvJqjlkT18xZAnCwrEVNlIOD4TWjOchYN0VKS7xMIxUZmkIhhl9Mrgb++DALOXBpzgosl
J7x87fAqhBaaSXIQnp8Wmbq2eXB0llVhESRdeMXjnYu0LWlypshlVD2tnUfi3fIuanOgfkUeggvY
unpaGulJetdB0Q69UoVHNGk7pQnDxR7HNhW4RjPepiZ0poefJ+qJ1/yFYiX8EnbPXVkZIjsb/aWc
7J2JiiVHbLgYmLLHI8D6vuAUOjsBu6yJ9UkVjOtlZMSuyLXlS/iMR2KWzAZi95DETZCnEk3I8Pq1
OBcz+8r3OHUOY1M77dxfCR2yUZKRQ97qCMTBTtmTt89Jvpsc+npfU/hV3msJEDKo2n5a9pLZNG/i
CH8mpP4AjET/WGe3DMOq6PXqz/vS9j163KbO77UGnO84crrS88r2dqkRNVKhGk128nH23DU6Vjm2
L3+cCAJZ4B4Gs5DzXRgyAtS+7CDlabgZRpvo3nDSlcTe0H8RBzlOYCaVUR//2j2bNgPPMjfKxCdY
p6Fz+IVshXoZ3P8WeYwbvkqmj1oEbHezJP1+df/kKRRHFQlMLKOqXzSY1aFIFfpxnb0jrPujRCqg
WjxyBb+WP8xkX5pEWf0MG8p+ieUZVCDNXlJQg0HH1OOBJ87G9wI759NjfjNQzuuxuR2z0EY7/G0r
jZEknkn3JlORmNZ+NMxtTLUF9cLLBoYj8SnAOktqZdoePyKhWhUyUild7nIL+b6yoYmKHPi2LnjD
vIBpPCMXcEn1anUEdmZzlL0lZ7iFqEYhdtMH2LYEA+AeUrd3i1iU34mXknSf/MxDJDNWHdwnrYGM
XvHP1/uVCDrBpGUwyEvQQjAYV3mkhDwEtfm5iX1zLoSOKQtvORm/x/x33DhNsCjDx/BEo+LTzO1W
4oTj4TJcBe60xRpTUhXDlB14g4ZbpbkyGVBGnTtdUuZHrneaVmb4k7pyr3r3TDzj8tNZd9hAbw3h
wZ3EuvUOHvmoEABu+P+nbHIkzQYbm/IJz4J5JzNC60os6rPAdppM9V0PJpK6mesUUjbQnOveVckR
LbSHJ0fMUVeqfjBjsIfl5sQamTEQEZC7miuj5KfanyOgSDlogS663/xJmNuQJBxbjzwT9moX9EeV
vgfoNhHXhhfvCwtOBJ+vu+vWJlrgp1ZQ3TqJYFFs7+qC1gAsHGeTvVmsv+TqzRJDpPUzLsHzXEyg
YvxE0SjSsmbZpRHzwKHDHqZMqKRjowPtN3CTfPdIQ9KIyXuQHa3G8tkpzkKf/xRP55NLWKM0dpsu
stRQIktu1zTrtca86GsC26FXfDdv3legqXcpjHRDYI/CL0bro8SqmpL2dLzIxJtD2bB/kH1Pc3yI
9toU3ZI9xiRHuk72zEnB+UIKAxgslphUfCPtEE3sn3LGz5/Urf6T+JVNucvlr8Zxc0cYQ0W2QzkU
YmAksevvXHLtBbDHJmnmVUSASCiwAx1LD1ShGpqD78xlUt+KqoHgU03nuSFsNqcE5wVbg6G0BRWz
BHhKIrcTk5N7EkFtd8JJ/MFL/2pBHK/7QrAHhRxuKKZggzmIxYftCA1JRQMYfCkKa5LT48Lbi+tS
X70WikG6sQPYkkI7ydhKalsCwtDXVpbyFlPY3Q8y2ELuguWWQtlRtGxV+V3Sc311efW1gBXVoyO5
o3B59Tu/ihOyu7V74Tca3RhCm6GtMQ8Xx38whWd7RQgQ+cHrEt8zyQrcZ3jUW4dqG7REjo80DvC4
gCO+H22vm69ftGBKHmMjVZAybC0AVqYnymjovko2C8mORyJ5fNyNxEJuuIaAA6AIgpG2ihhCXi/k
SaVaol/KkBuroa9w10RTV98RUSSkUq8yb4Wgoo01KTxG6+LJ4wzn/VDjHJdCSzeTgPsz91+iTXrU
ASkSlNh8U3TFi5jekaHdk0vV47DiSIlSIpY7AbgD2u8RSm4UnVjBoOCap3ldWjZhLrsK3yEh/PSm
klEG4sd3nSet1F6HuL1oWCSMI0eGS/MfaKjr0OlIS6ncNMi/ObtO2Exb0Z+VDWO7QpUH6/igpLuC
ikL51WM8TBrAzqOYTvKEN6bX1W9eo+P9MaTEIfjCVIUTFhLN4cDG6lBdCbMqmwjFMA2Q7OxrvKNY
BOzpPE0ohw9irJBY5Gl6cf0AJH8ieN0PpucWCunFEJ60XMcc/4DD63aB0Vrj2UdMkcprsoJDwa2Z
voA8MJgtZRb7s63iwk7pepYNTBHe9kzQQdLZFaoBNUDeeiPebO61R+u3VEQKPmdofflCBNQpC6kU
qOa+J5/AzvyXiCAl0c6mrxVJFloUJPHKYyW1yWH25Oygwq0eGjlBBWIIunk9vUYR9V8i2vezKpUM
glJsaGREhsMwyAwziPIA6/IfnrfxJjk80n2XNIJEbgYK/VhZDBc3dLmFFWBJ9Uq8JUbmgA0Pu0aN
5FMbW5y34BX0o34z+yDHsw+Nm26xJujjPJ6Ex+Gu1WaOm0AXLApaHT9R09hZcrB3E821pnR8P+mU
EiGz8VyZ2IzQ0dUAMDXDwVrcMdOlhw/0vOmmwdC7wV0SC7LRXnXLjutXFrp8Km4sU7nAc/0rVoVa
xuaTt9IDY6WJEomiRaucgslkw7iWwTfm7pQIzIYexncZYApIQG4+dNiq4jJZIL+VrfSBHdA/53p9
Qj0aCuJDtoSi7NKEqbWkIY/5vk2TDWDlgtbp8v/l0+oksGgw57Scn+uFFBKMb+RjCBiONhew0el5
Kh/BQunlznOycu5CcLqDPUn0uwHQWYEzRZHVzA+3CUtohZzwN1WzvHekowN3DERwsQoe9nidnMM3
5YqirG8KDvnbpupzb7/J3fena9OBu3+YMZJDqA+2v0O29jLuwZVNEhp4lDfsj5W/ubhF7BrLh0x+
8xP52FaYeF8zCkeaLGthL9cfNouluAak7pre7fxsmHsBHOCBjiKgruk9JGzpxZcqKfq+CrMZLhqd
R7e6dIAMXLOZ28JLFGWW1QYaw6iaX/+OrAKLyFTMwlZ6ALDkx8XXUK8aOMXkXRBq03fsg36tpNXT
Lic/7x1a1SYnhN9OVTwyvhG3xId6T/Glr+mJeAMpn/ObSMYYeYYJIpYUidhom/hFn+Yfl1UyDeNm
6etRfixlN7BUgPAvcDjuxbgucGR7wAXQAbbq8Ci7G99u2VNWR8o0tjK2G/FxKAEQcjjwaojFuK2P
h6LBrNJJ/SF8tmNBqfYEFHDFCxGfBpD+XC9xqPggg45ttIhR+PP+svz/EmAOYj+6hUP4xhbF1Mfi
gifpyvo75uJPalCJ9k/aYFvNyniZV/9sNqv9MBl+kyJz2JNpb64tPSFt4yZo+c83dyIHkot4xX0x
S9CL3+RLzKRPQytMVcx6dCQjbOo3iSx+AH6XfewEObWKlGk640LcfvvFGBw1dABO7P8YPq2+TC2P
k+CIn0cWfHCyTca27oXGzGJdUdg2HN6p6C2AbJParYOZr+yxCbZzqvc+xJvifwgIuDrHdofp3G7N
81kBtINp+AOvV+Y4J/Z1LFxKKKDK32AmFGCS7jzKWDYL+V85mAMiuXhs412UWD3Q4ZQCGdUE/k4Y
8f/3/3DksY1B/vRGoNaEcGAvyFV2cAH5XTCWdETxkCfPiLnspRgGxzZZRQiDyyv0fT4yXTdC77yg
/0LDnQPyplwHBeGFGynxmTsUfdMkRqdSD/gf76l6zyJN5XQFQvzqzv+We/jPz8AYWTYZLQ7OfPt2
c/gcomP6d186mrVcLbDeVS5hji88RFIwST+Sb96ZsmL9YtNvURr443+NMgTCilfsxitbgggBxuCV
VxTA7tuJL3NQNKr1YzWmprsafZOF7tRaQWRb/tCbWF7WsXJXG5uNHGuBmDhgj84Tro6jKr6cOG+l
VBq8ENsw6wxFK65/8NoHumUs5zRP1iYLBUyKJvQAFWKQR3yLv0NGu/6fI4ZlqGL5EHp5uTv2WMXl
oPalwYan5HBd3TZqkZIEWBR5wthiY2YCuGUK1OJqMPCbMzKpbGscQl2+2073vaeV3zfldoUmpjuV
tpUTcT7Ogc/eciPA55mXw0a6cfAgat6hTh97PgLvT68azrAiFSFdw1EGTCg0PfCVVuurp7IC0M7h
WHzkq8+PQVZW+PFecnrwCs29tdjde0uVu+UQ0RdkImnZylmsp69MuLXMk/OIpfaLo8icpSuOB9MJ
5n6/dSo+8aQ06ExHjemGQJYtbmd790yY6nhuTnuhn17P4wzPWqQv2mTEhcaZeyJVKiS0uwY9p91I
X8qcl4nQZXCm3bTYQVyP6RHKip9yaPjt637TfK/k5crvfWGvOrlbzKl3t0VeraP7tTwJmVZRk/Qw
61WdcWRqskuERHbxc5HZFwfj7q7fc9cvYoT7/iDHHanAcTUR+x1J5DYX7e1+rrtO5v3M0w7yGnmU
qNH+P1nHQ7GuWTianTWgKWyh43zX/E9EdyM07VlhN3+9vO1fy+vJ2wpMr2lRw8BjFNWiz51e7/uR
Mwu9WF/OAyO0NMWONZq0vOxR2wKOcoaIgtTDohTngjPLCWH0/BJCb8fByYhqTeDTyxmKTyXW9tib
5gAJb1IVzC58KMj8534GuUdKLHtlJz5DMBZnJEM9EFSP9z8StxIXSM855RwMUzYyqoSI1Ovyp4Gd
QLK1eFniho0CB550qM4qoHIzKlbvum9p1m5CKsckDYDrWzhJ/ogp/bsgDPXQIXqgUJPr89Lc5m6X
BjYeiJ0SrieWFQj+hh2kClOX8W+PjkQ5NlXRVtVN7g+NN/6z10zJfN5wSQbGCJPzZ/xeu+jLmsud
Yv87+gtilTp1QH24Q9Dhn2JdyIPw90gqwcb23RgyrRlQxpqiz+reHL0X1fS5m4vdAoJBsZygiUk1
1XNsvkRjEHuUBLremHltg6XcwBo4jM999iS45ut8QzXyeAsLtdw+p3g8LxOXLaNE89D5xosP8B2+
yBTklsbadi/HebcM1bNOhbG0J0p5zqSzRbdYVgS6dd5yZ9iB1iYzZ5x6X23qIY1JPnHQmIXWCdUp
ifmkra+/7NDUvHhar39x9oF+fq9DJ8+1P0lfogiuDn9lJiCJQth3BVZlMgmyEvy8Wwj6oVFE2rGt
n+lCtJkSvE3RJCo/DjX5ETOpVi7nJLDmQLqE61yN5iaEJSUIOlcTbMfL5c7B5kIdW5csmhoBlJrS
ePBb1sBROzgMeuSA9rGatdQe4mCpaUMe0JwCU5M4x8opNhLnAspQE0bmMf9igFfexc20S+5XYxWS
AIDqns2cbrVCzPcot3fpG/UzLit+uze3W6KFcHuqYePHUBdzxlR1fpnF13y++5ahUDVBocIiZnbU
8cWMuBP2uF8+vLzxuvbs8B2/taWFMF4H8VuNhA5tlCs8qfcXXV1FWiiJJ4CbTIQoouCj1CcCMBu5
hZQax8UbIFqJBgOgS/7+UoNxwsL+kPwEHJmRp621HNjDABpvnM13z8m1ACFxbqpvGeVJ9/RVgkRL
mBKlvwmUpXr2ThadLM3QmGuSS9UHTpGe3ZhsCgXcIGW+YhYi4YfdzdnF6GlV/FbcugB6jr4xuMs0
KOXu6NZteS3Rm1dGb3dNiopVCDGKBA9nlFBcvJAqdBjUEsVFW6jVFNoUH0R1pEBo1WtqWnXtVu+W
eWrjrBgcZe17lm5GPo55sqRDDqV5m+d4zNhDsVII/bDZoyjF+XiTNuV8bVL8gBFnqj5ARFXIcayD
OBOgC2ALGhDXEcttewU4FudUYcS9uYTuiUw+L6CoKAR8iQlILsBc/YtmH0ksGNszxKwxEejUuXD0
J8jYRXOb4p4iZGZITUpyNM6WSrVkug4lt1SGorNaoWNu8HNv40G5mJpaXPyc1HrTHC0n4CDeINL9
S0fKYi0mN47hgqaJeLagAdM2Sm8fK83XfY22h8qMtKG6pBpZHCvxLjBGmooTeCwm63bfWHeCopjO
dnsU8XCeBOllO9UBBp0aZArQen4SnjkddpkcayhnfPsgWJ/xrbPB+SpYYbw90R+w6YBOoIN3y2D8
c4IA7SQwtb9pIO/lpdCU75eIM6u9HccvnNer1HAVFCb46uYOMjM6O3O1Ko3S7hrB3NLZRkcCbBH9
w7wHIvIXGQ5aj2H+ykmVIrx6kHWQ+iukGH8nI1/wVV+PX92PtRxpqqx8SBGYxlcvCv4TyJuXT+pP
M7lA9ZuVCF439mnWhOr0kR0Mh+02mp/65QFwXNRnMRsQTnHTFwo+tN2OK0CPP3hPLWM26e1tLaKw
cAGbsEetN4yHHbEXcxTg3T9n7o1LLHjosyKEwKJcMQv3ho3WnvQk9sgkowa6AjnsVuSWKz2r0pxA
nS34Siem4tTJJdgseJS8evPPv3Ma13oJPfnWnp16Ku5dT8tc83McftGY3NV9qCvGXhMIfPy6ag0K
pFA0b1k9ndTp41Nmw3au2R0jE9Afp88FBjIK4udMRzR5xU+H9gC2XxIKlgSYbveKkyoTvfdOTFTY
JFuZi7cInljXCkZTjB/RT0PQNEGzll5FYC0GRuvKbUcCnAlkltby+TZgY5KrKaiQ3ob8BiOjnwTX
sk/u5vyWVG/ECUpuLU2qbkGx3ESjQDDWyqCs7Wzox6WCXfFa8ny5EIsL6qm5PiuPfemvF0CryCKh
HLAqI5kqodBvZdsiqgjJ1sccxoRyLuRmzKXTNCgvvx5II6Eq7DQhoKnxnfXAyg0YFfDUT2hXf+qR
k4E/OA9Xq+ShLkW02TAl+8PolH8tyTv8APR8kFMD2sSCV8mAVZrVb9tIBDjtl2vvWwXLKecylfAX
uAO4BQTKpIcqSvlEQv911N7TI3wNhR2dn2s7rkfVW+8xGv74p0PB0JjAyRmOjkI1ir+DgfwCiUqU
guZmwPl3irEOIk+fQArsFJcsIM5ncasa5SGM9ihqKZmEo0fArvCPYQ6LNwZ843RTxwDq3jqwl4GB
v99EVx9w546Y3Gww5GRtKGBAxupAuQbwwdjsj8Fl+g8emEWNsJdImlQNJx5WzbR12CE8vJlKUlo9
I3EREDGkqS4Es6/oVZTpveJzFt7yHVAF5tADznyzXUyXtJWJDrzlWqWqfIcGJNWAIqkQMAsQof+R
v5hlzE7JoVEoyHRGm3EPxvvkiWod4ySVgQYoZfQXokmTs4clEFyzCTVonlvuK31xqrJyGQIJloHu
/Fc4JpMrUAiD0OB9J3VcKdJSE4Z+BhpFssQayaUA0woNi4B+l0BKqD1XNl/0MhODX5aSL7ws6iI+
tWrE5B5/Xy7PlKbtLgmYrPLvbm+jBpiqN04z3M+l7QXmtiDkqt5PyUr1i9lRJJba2yohvl5yMs0K
f2Rvn2vsOhbDS+GRh64MmhGIQTZeEyC58iRbS4B1B6H+KlpkiOXAoXvny9w4NzlR2QzhzDiC4SHe
mKIBKIROrcY/vRPNPKx7aPiW5HTOMTBiL4XXedtCqRe61REOlJsqwQWa7dFqpThBJBvG46HSpuaS
3fZZGJSLdcsH+VlRFqlRWwt2gsq8ytJQ+kSlE1PrxcDHW2Im+Ge5pEp1tt3yNRHzO9FGm4a4oEa6
Z2OvEZubIWx49Uw/6aMU+89P3pReuAiNlF21N+WA+BWAA0NViY/3/uSd7/QYuXRBoig3F0clpCYF
br9Yrg2k268guyemJhz6OUSJE84L9Kt7L9W0lJqi4xOCKvx+sq2ok+clfdeIAFpx75CHOH+akPzj
u5ItZzS59jdR5i9uOKI/l+HcZK6XabIHcpainlTcgKqklt69A1BvoekExvqc6B2MvHiSksEqgihJ
tsWmWbJxB3LvKfWDWkOYoR2D3tlwdBXDCyIcbByKS9HNkN4hbkGd/tkXe4jTBh8V+z+LzXdJ+8mV
nTawinkww/47gXGgVrxPdiQtXD5n1MiKLk0bgKBOjvTPDf+aJRC0QOIRxo58mD3o5mN+ICFgsbov
8jh7xbJd0kczzysIIO2vra3YeE1KhAPMa96tENXoICDbzKM4UqtDnbhodEo1fi2XODUR44dGm8nP
isGz+O3srWzhzrNH2DZM3R6HmhoGVcL9ZR0OJ+8gqGUqQ7M33AHALZoEjLTM9jEpTCCqGW66Ovbh
aqyN/hesXCI/Ep9gwyVshwf0Dbth4a8I+BPDPQ8nLQsH59oQOwem8PJDfzuxktxerBfVEw1F4Ryx
Lqp/k80at9n1/c1Z6On7fVcqq11CONzWaEi1fDS0GR7UCoDpEqG8faWNnXK1bc9JSOHB7RQOSLum
ISp9MQyxyBxHXk89DWo45BTuMmGL9lf20C5Emy4hkfxO7z+4QIGdJqugLUtGWx6AuCL0q35eGl9R
YCF77jHUZfQFLuVzF+Rd6xGB4ROX8Oeeg9EpcO1lUSqxoJO/Fp2DqNWm53Os5ZvY7CZ6z+/+iTLi
/UDrvs9ntdUn6EmLZE30CFglnIQNbX81UPVpgqq0Ue3oOaz1AtTdb4TFMZ6M2F22nyomQQ/WleuI
KN0zE/C2KabpST1BPxvIBWdZIG/wWqfOXaJY8/I1G/pzZBcFq/wafwlROpHv6PcqLMUGMkZgqPVU
gwRDYzdvHxIypAPc8tOxPzv2hmHTUUvziND6iUP+w6x4567a4FKF0MPyZ9ZFPVoUNXRwvHeNN8vl
c5plRAJp0+W/uur5QTzrqPpMgO87SJFAavJKJN1VZ04O09lCyFVl+eznwgy1OhQeHSG+kjHdoDfS
/51wqDHD7+Zh0n6ANTAcfXn67v7lQJjsqZAV2KLUxcyfYT9qCJg0/dK6lL+rs+N1cKSdO0X4F+p+
BfyHAytOvdibSUpwnDz+hB8ymBEJ3Q2hojG8V95bnvW6N/WIZEdQTqkcHE3FCFYrpGurIdqnTPtd
/BXpfnQiiusou0T65NnT24hIUgU4jrXtFZhGJCumDD6DdJzpZmoxfAvPuHnXBQZ4dJ8Fo9Cpqe22
mLk1kNIpdiUxdCdaVFYccV4WoPiylJ2lOM71PT+JF3jq7WuH+odK+KVS3XCTdBy9mvx1MpZ7NR7v
9yrYDGdHujIKZT05DZbInLze0AKUiNkQh0JEnrxKLOSfiT5jSXrgLe4yyk2eENphilYpr019YVtc
D2iwEaTyd6wDKFRi+T7Qw7S5Hqbi2PAASRMM2aXXIzQFhDlrK3PsjYizOLcv0qSpB1PtXDh7c99c
J7HshQMde47jAJ5NZ0YvTeO53GQcPKlszWDZZobkn8LjCmK/ZVLNtr2WRDUjY9qxqONdiOqZhhfr
8wnqOx3ieLTwiInVmRUXvb9iZNsCcw81tAjEbJMg6H/KddQglkzsK5m5wOQW5CkcbOk0nYGRKY1h
l1gu1VAiyJhbLCKm0OjTAcp10UUN+kAXLT96smjO9aPkyy07jRZHNk4NpD/6Ua9yTkUPw06HIfmq
ccOenD7DdetgvJoKFgOeRLZC3iSTdIZU3WRJiveP/7c3HohQbI+nGAi4za/N5UJ29HQvhLRHPaDB
oQmBUi4lDGrJc2z7TeAL7cFw2ZWYEdtWODt3caacnSbowZ5vLrvIc50wGV1foARsUlN/OnPtgUEN
A4AWazIDrMNuZXHpGGTGsK2IlmsLvvDYNl5SToTChS8jx3ztOnioZZaL1nCFmHBCdMOfoQXWIXEZ
FkTLKCBW1KhK+lPSfWMHeW/l/Gl7VQ3/A8xu6PvOrw+TY9FkpyrPpYLiOV3Nyp2GUXyDbgLNrrTT
sRSCeiPtJ95Fca1wUvYY3dCvtGASAe1W5qC5QwFDu0zvDDo38lxdURjbiL8foIY848Kb5GlNuoPj
B9/oO66Og6aPJLfYYMVjDXqCM8uHJRbmNHwFBVWtPLzvKtjz3VKWdMlm/8n8tq+NxVip+5qbBgu4
tUfTCa1XOvmNb7aleIjkXxIAo3wL3WyDFsJ6BgrKtFDbJPiv+IQOWes0yuPEb98Frn0Qdg2nf7Mu
ER8IDGCqmfnPgFl8qd7XblizhYRuukjmuakMXrQFIp2CZRv+bzIZ0v23MmUf/ics11KMZcOGkxA8
LeceJuEMNKMNEam8upW206LwQrpASYyW1QHjqfPIDWsgU+UNPqM1cRW4KqzSMWobi6XhRUs6fMWR
5UZbUX2N/ByHYTPMV5WVf1oMTBrk9uouGVFhCRsWaFf1CRhNE6FICo4nWSN2QkWrzV6l0FCTJ9uX
M58hsbtdF6PSw4MCud9jvg56sRiN+dzAbC8SxseeEXyNldIDBFA0M0UHM8u6xMB31kwYusIJE/42
bQ+uh4xjJNbDANxIEosxVJaMVGjfJFlY3u0IX8K/mq4b7zyPVswBqkHxCwJ9oBf+7mnVWMvsRTM5
sjNIT8ifynZAJc4uUdSDlSZy+jKqju5bPvLj70sbk5ycQR1wVtpr3tv4Y+DkSjCdkkQrZ3yzfpM6
Q8iRZxKWaxF7F2vwGh+Al4viw+wiY3DeyEeuDu6eCEXPYN8W8tz3kdrVIfbrdmGKX1nLhXgltHC8
udMLUcuaOTbo9lRAbM1fX/CIP56uVRD8g5LYxRyzUIjMAxeKux6d0R2/IZOU/ROr8D8WkG1KQBIq
RrmP+dfDbt48RN+38dULaxAjds5ES3OZrJ9BfVhQJNCkibKSQh1GlQcY/yErz8m0HEmn/ou9EEqC
qYV0AZHpl8DfluESKYf0ByZhQs1zwXKzpucXrmlrTRzWRYKK8sbDO9HDGN9iBX3ki4djjG6GqNuB
/SYn6u7Re4o3X1IOPotBnaGcwfjvQRvR0GvKq+pVoy4rL8ZmiInNqle1f++2lHXT3I91OohcYa8W
1w0f7qGPxFktNl+p8UCjg+g0G3cZhXXQ7b+I2YbHbPgJl3JXziXhQHtqUVlh5URum850aFrS5h2w
bIrv0bhEfDOQ/p0hr+a0vlTnuwDvqf+Ck0EIaixgcldzmnDNZ+BizLRpLJUDoltolX9DB4XIXQx3
+SRbeWIevMCPMJFLdiuq0DLdEiz2llnSTgM/eQ06NkjMOr4rYDhi9dhAKIGhynhWeJJAw3IcCn41
GAMhxMuny+PG0oh81hy//HrnxDFUyrXyKXSuibKNEEvl4SNer7ydvlYNrE2w9qd5sRe+pxs856ca
c8dm4Ljr1OnmqlvLjVg9JAJDFsmTYGuPcFuRcgNUR620EzvHjEcU0EekizNIQa0fRQrqutQG5WvE
lNKKaAwUYlQKzQNSCIV9nsrNLV7D59drm3PmkmHQOfh3T8+h6JyONBG4vZ4jfrgleNy/zfbDZIav
BZGWIoUjyermer4g8b/N0wMhZYG4S8w4Tooq1eM515V4oUxm8AA5w0DbtSIGVROcOJJtCOljmS4I
JKTk6t6Ko91MmWNsMtWYHtExZew2x2+w+vgRaEP6VHSOxjr0UtQfty2oZrqP1Cs3cXxCaqaPJ4tF
bhwv+YQA89to2zMmNOQPAdGzjwWr+DzeOcpRuZifbtg8/tbP+pG35sS789OrS/a5PyWa+VCowV4d
hzZZWdyEtE7ZdRqGqbcNHFb/boMr3K0ooa89XytB8eP8vIk0LYr5vsmYLTujV8qt30seLpQ8Sm9a
J2dfZMI4v/yj8dQLoyRYf6n6/7YRZHQRHWlbElbrt83/U7NZfK1tA4y8UCu4J31aVFTbzohaL/oA
+qd/Tf4iv863XP22u1CHfbsVGIVW6c557cWZ7+N37LfT3drTDGwhJtSuGYhxyfKZbtBSIEZfw8xQ
8BOsvEtEWEOfnDGTwV4UUPM7h5ygEaiW0AHSLSmdERKK0upAWD7kIAhdW0endpY71zFm/+j0zxHD
A6KzdQorR+d44fjcbxWCpOAPSgxIJwy8ehnZ1Fdpbr2kKMOfff0CTg3adTeN+aEpSgvBD23iF3EF
MNGsZmxNW/tIVRVDt3RdfKWYwfJmwHeyQ3VRAwyUujWUMxg3LXHAqSsFzkdpyimEtOWB5QSPcK4r
6oB8Toh31+K+ZrXhU0B9kwwwaDxGzw5fIBW/OuGckFgcrxPbpU9IYXFFkwcDTvzkpt4/I1FrW7R2
u2r43qo84wu5Ftv33egZD9RL9SMR0F2cGlRCh4Xlc3zMcbrwbW3G/hGNeb+QJ+blWOzShNLoFBdj
KvQGYKqX6/foKZ0WbcvfobPhWrh0YGLkkJ2fqyKjOAfdlC3Sbggk4ZidFedgpUvQpFPWVcEnefrg
vwpNM/sAZTEJ7v2rlosNtWDGScVM0v8q5UDvwdOX0xg2k7OAh5GGrZsBJ8mMDaEKGFJTzy4E1njc
SnE6f3qygEHJD99NwhoiuT9znT+QXV53P0Hmejuiwx0ix8HWFgCO9FTLot6edjm77jTUqG84emb/
sAeK8tEgOPCychsPgA+o+3N70M+1HuqI0OK7qcFo68t14nhMvIDZbNQVsZn45Cy0+midIYGurZWv
iB1At/yTdcLMJ8gRi+/64KG4/fEvTtc0cEH4v/80IGfj/yAuW8o85JFPGiA3tjGbTZCIaySecGM1
UxkmEuDvTb7S79X+X0h0zCgJdzKxBWbOX79EjhdBh+/ZfG+0EO0331V8gZpVojnLpbWmEHSg9UtN
FqYs9pUIoCJfw4aWhlK3jnLmpi8OSMJR7VAh5nmyyuTidga4nJAnevrYDhsvS6ruI3bju5f08W33
Lk6gVy7oVKYfekzpwkzSbPZ1gcfqnwdULPN9K2c/onBnexPYblOBecL6muMSyyg2lRQkX/XJs2jl
UiI1crOWN/Oou0jipSqnlHDZDTEKfWAjPBLBY0SRfo08ail+SXkhWnJIAL5Fu576iTNr+l2JUssW
3LYu0M5qcpn93L0qAk5Ez60x10vtKm3LBYUJGaypUFf8q52ST15N0RFWIL9kpeQDcB0EPT8xPs+W
96LtqIYKUocx1lrmY+dHnSMKJAECORkyDbSZGOlUEieqAxjMmLep/ocoWd1RO/Y8iVA3oCmTR8Ve
4XNeWvK8udHUloznT28uRlMxJRGKkDb3SdkjC2oIHvkpLPa8O5OjSPfHvS7zw0ghT5/r+6s+XS3H
ZzoBxv3jDa6kC9dBDug/nV0xes9TfnpDGXIbyGanhpvJ4/5oR0J6BKferhoUhL525HEiUd63+WMU
C9DlgGRjpmPQAAx/E8pW6rO85JYXCLPaucuwRUYTXwBDgDxVtapon4at4MRoRnSJpWe0Cir767s6
cRhle5iNr6Ho5VDWs38LvGgshvXEu3uPcdDPatZsnoC1nnanhmim52pS5RepeTAlMIFhZMRrc5/C
fa/hPakDHe83InMtqII6vKNs7BXOyF7bYxyTUNGHD93Wh/YPZiehcK1abZ3Ii/SNBOqPmgaHl9AR
Nz2E6SH1yJsbEZToiHl5xtlkA8/dLf5QfTNJJIoL2VMigUfazFjgKiga1QxSqU4pSNy5BFmM2221
Qm57zpUlmj2PFLRHK/85Kxm90eztvAXMMUUL7LytudXgoVgnumtJ6OO0FdIRpaU9k8MkFPcJCKmo
pjp/mFn4qwGibxn/xy3g2tXbaiKvHUKiuuceum57Ctncez3nAzMDh3xA9QFU0L5Y7PNU269PKuLh
vUGwpbey5PekWxVSUky90sbmIOOomUYCp0NnP9ITZPD9DXIsoYJG+LzjBookie/GxnjfYTKO3fEg
+gFibbtco3hAMuE7nOtP7mVlhhloTGbsWGiqDwiV3xCUp3jzXhe+wcDiVI9FIOsPSimI/DlqszJs
RkHudSQv31g2SoYO22d3vyP9RuT+HS8HrdYhTF0VYudZpnbr3uRl4LGPcHAJModhlPtXffm6Ayn5
Rvvhm0Rq8Aj+AKmnayA89LkX5bEeQsIt/RvK730fpHhpTXjF07zPqysLdOGCCODtx1a74xLeGco2
ULmIWTj41nwS4bu7iPYzKsICXO5jMpVd3IlCUhfQKqWPa1qMhhvZ09cGqo1POk6TVeL16oW4H7rb
C6bU62d5TEtL0yg2aPqDpiQL+qn8vbdNteFfh7YlW5MW2aoOG622Llb71n5mqm0XybJXOUoyyr3V
O0La48eR3klgYSKo9sGuKJbX7EuD6riNAdjAKdCCV5FiTN1PXlpZYSO6by6Mn5pohDlWR41VQbv8
/ZeO3dB+dBlX1ZBZ8TdiFXwRxYxyQbAIeODtqZhwc4VealCvLgyDDEIMjMxJqMa7wt3uZCmGxATE
2och5b+dSvigWpw8iKdr8NXR+SxkgGJxLEqVncfKzk4iBKWjwwA5/M6dZ98HTpysJbrxUONX6VXO
NInvOjKWi72teWBiIOFIOF/DAFh9fD6/NSsaqETezalDdqKbxo4cr1s0DUho3oEnwShaIzH6+2Vj
PBnyYvRvHlqeS1RpxpB4hRlb35CAEn70yY3MfPoeG57ChfhjLQOMT1sQEkO4fXnnqElJtkaBuDby
Bt8fvrJUJAtp3Z26751BBUTaXTS5EThbJ4OiSfvr1H7vMw23Zt/EKTgwPb9rTfR6deYPaggBOqoZ
TmnuKj8iqxrBohBRwXbgZBHhz6nVIghsRHfk0I7wVFMnFO4sOlMIZFsULtzFA7tz4Jp++5q1EEKJ
eyhQmnwk4nM5yxdbDbUgD3+V1ML6tF2d1bqLtvQ3q+FmeQvG/KhTSJZJRlSrozax54BN8fUnk45P
8ZWkr+5v0z61y1t8QW8/KOsRTkko/5YkdnhWrCrztY11iGXaYmsYgSGdqOrl9zXU7yvdiHrjg+37
kNuKMpNK73c1PsJ2NjnLY46WzJUDslut5lWNLaM2BwvvyDtPrpDpN7XYwu4lhISqADyrHmiSJXKa
pOa69hB41hiqZUcp/1INBmwdrDv9w4TgXBlaqABItWRMOQZyyIsc86yonZ8cb56tyDby/pk4AddT
h1n9zTRaSKk/YRYydEpIn2txplMkrd4lHt+1VB1CH7DJ+Mcv1KhxgsVwdAsy9dco+gFlSyCJ2SiX
ZMJqKMseCpmLSYjiuawjWiWgu1WuIy8xelMACY1KzzWevODxYziV1BE29sOYIWkcrAzKCuyPFoQs
oim3E029bwpFuFlJYAxRCeeWzDQJO2vrdvuURxysIL2qt1CHlJRKKOW6xN9NKUa13/NO2EFMIruB
idtAfnk8VDgNE/IBGLBUgWatmd0E1/kSnwPmSi+VhVhdPdm+t3InIg1hrNVZMMOgWQCAoUhIIxB6
ZoC7sTWetg+Sn5CXI5pvhuBBMQeZejDqCuwRxJ2DuWQV15X/tHECj3Yv0NJUcHqmvnnWtm5VN110
dsXDsKkP+iZFjCD3bCLoxjHIcfdwNMH9GPZImHqP2/TFr9zXrEf6fFhERqibJ/cgYuJR3mvDko+5
TsI2SOEcF4EwsRaraw9etBN4W5jOkMseG/TP6Wy+HlcBNjROacwArYhlQISf0Zg+lmZbI8TrbJPn
BRMSzuIzQRVV0QSZ0sDgXwyHL5D4TXKkMpiNBgS9d1jCFgMN0tESLku7s54wOObAKfbgL8pgjcnh
SBtkBFH+Q+MSaujs0vj7WVNQcBXb9QiPc+fkTahMHi16kHcNnfxQlwS2FsBuEVO9BIQZ+QICzqOp
FB+SpnaFz10ciGdbWzNYc4A0EtzYXBF35o3niScRPLcjS7twUMwR+dSUbzH8zkGy5phCSV9SxDwc
gu3wrLOWyzAbC3QNbZBT90AnfU2WjfaJXjFq2kqALlDK0IdVRkpYum/j/NsnrbO1DT+Nqw8St+7b
Fh4g1Snca1yxJZUH1xFY/7q2c4WFSkhRrNmKK3PP0OL5HiEVuHksezOZ1z35jGzvRvN0x/7NyPIF
7zWVs9LUau9DFfs++0l+Fi6vDp4ttCE/symaub1rENCmWCYp/4gkzMZHs14rcoC9/u7axFw9rOE7
IgnQ0rmD15M0S1YvreaITkjG1HsMtjIRAusGyx2LRIsbu3etQ+UryccpU6ALfB6lb2RmIWhMk6Ak
bGbosluws2pJRzjzciWGmNvqfEsuKsE3yu06bmso+f/ngH6DOmiy4gZspYKuHUxcSjtm99Q+52ts
SUQVVG0HgxrMU6YJRROJ+rIUr2yO5y2o4YlNZPYN1vbPtkYM2DY/ioxTLWwX+cvnSdwZWazVl46f
i0iUng1SApiqBtOxo+lQUlpjOdo6Fc/dyP0vh86YOBphmqyxI6mHHqIksdB03bzzJwVq+ZEVY6tX
EweV9ZUoPY4TZ0iw52dZdsfP9ReHRzlBfQFYsT01O3gT+9Pi8B6R8zQmFL9hnfHWElTuZhNAdYTH
EM7eMIPE32Ixs6FPL4rHN9ZSVN1BhRTcg2YANDv7ng12QkDTwemChmSrYtxNc6oFbWrcBd2mVkr3
3HJZ1xqIFXYTxX0rM6JYfTOAx5/8uqUCZk2VS9fuqwKUhgMtc8N7KduQcWTxcLl+X4HsOgWhgbzt
6qmOnsvJ5AyyZwkVPEETJYreqfky3skBqO7Sra31kHQ8qur8hV9N2LsR9giCoEsTx8530fzH7YXm
/XgXAsvy0U1iAE67CMXT3NkSlXD2H5leC38FHmLVR2d+sLMtxjzUa8X/hWuDe7BwgbBFn2qVLT8y
4IfDqn063wC0tUqBrT9Z8X9rHzvr75FGHu4YfSrdYhLBwdTpsP9lc82HbwejgfDUgIvos00Ww7eu
HQb8GSdewWn97OjMBybpiATrioKOokleTaCAUMIV5bxWxlTsBFsUbrBLe2AHTBDo/v1t41EOgE1b
WJuk6dEXKBa+kQgDlbMYnMItCEP6/t26iSV/V/rWv7PRqM1TAFaFFSOGKB6Gr9p5i9SMhkEZkT0B
TwYt+NJDWvAmrpGDRbh1pXY6KDMjWZYRseZxr8IAc70GujF/GdhbMFwe22WiwBhRDSlnQjmEA/sJ
Mutxs8wTBRvbISPzCWuEj3a5wlaBMJ4wPF4HpBAOvwSTawxuaNJnvarFEros4ssBQUGnWbFi3BBV
Go6ATDdeaS7eeAZ9wdendvguopg4hOIJh8akI0mLdGeEzhL8V7V8WgdoTaPSsiU8hIbph2OQ/cea
LYic2CT3NPz/lzX0rT4F2JFb04oVli4cqYj1pq2cJnMl17Je2bmVq7oXCkAzMxSsP9yeTQ4B3of+
UnOp1wcwg65aAndUdMn1V4puIxqvH98mY8ojc6yrjsh+wdTZggEOEbdseJCE+u6Rsh9xp2i3O+Dw
v4E17NiatIL9trpA3u/1uyWmBpTmc6JpTKgoMIWYgkY0g3irpGpyT/LV9WMtbsm8zvpCYIGUh+rM
qUM9HEAFFeBqXvKCv2mj704aRbc1Pu70kKgd+MaFiHwbdNq3yn+zWOkwtbeX9UZHiE9bKgryrPF+
uy53lK8kaA7IVinLH3z8OJzyoU8vJ0CHqVeH8LtDUk/FVaH+4FMIJcQW5h1Jlr4YxzeriJjGt1NE
2NOvd25lQ5/4lprGuUPc63vYT4RSvEnwdKOo5Utcwe6/i+VmSeoGr2BKuh2X9yUb3PVu4nq6iYB8
2tI9MyVhWsgS4wWjzQdr+79Jmi2ALv1EAuBRZUYIPBqz2GnO9ByL2Ntny75rVRtTnBuaw/WDE0Kn
CpddTGPJjjgjk3cfdw1MZANsqruiSs3laW+d3Zy+Vd4jn8yBg0rBqAniIxk3NK4QdHy5MMLMm4J7
sltEpYKGyMI2J2iwWpdNBO4m25ADrhkni2zQ/n5KIcy6qJPk4K3FM5wwA9xYfQwXzX2SHLCWmQjr
l5qHI4cEl6qeF7/i+nEwEdOrjShexhU3oN57SXw5HGe5shT5ik7GRKMfRnkURag3dgFPBUwtmhFu
P/BpaliWWaWkGIDtPHC3JwwuJnm7bQe013p1Z8pwhyFlwbODq7wb31yFxVz7eOqm4QkhmDFv4gd4
iqLx1+r+BawJCx0lJKByutZs01rwR1eH59HMEQh0ermQWwZDUanjaZP8lOhV7Ne+Y/DyUPXnCbQr
YUcMwFCUDRMzBAGtHLHRkQeRxdB6mzV8WFfZKSeqSzBi5Q6AooIGa/4rA67EV2t1QHmZeJ7Qw/1K
g9+KwPbA0L+aGCP0CRYbyI0swWtCl4/lGeBlgvjKUbUysYYfdbKzDQ8Bd/9wGs/fPHuvkPOY9A81
jbM0vNq+JqPFwPrFz9D2cgKdBUkjdcKl93Zc+ofJD4FgolErnSsK1RIjydb2zoJO0O3yz37pyTYW
55ByPnB+8LTkpwDQ2qR9APL2K0ZL/9MY2FWnms1/R/ffru2IR6DU4s73+6c0DkcL6lD81hU0zsJW
F9WrQYR3cYC1oqTq5GIqF+fM7BRSZwbPZdMtTSBHOcVeWUkB52HNUqhKKBluau5MaPwMp2O62/lj
sno+2LNDxyDuoaM5ULSHrXX2E2gNGql/wqecUuGFzqHxfFC2DjImljsBgQOTfiZadHhP8KUpL9Io
KoRShWF3m31qt6F7va2z6FmXtgq+F9z4HAjIzAICx07gf707kjwrNKFhw3BlHSwsObOU6Ly2qxzd
pvql2hUk4w2wL7UOSf8dmqRM9JSfV+zEYzfTNECBFObXss3sUtt69IPEOE7GJ3QkqmCK2vIQKp75
gIzxdm4Qe8JxO0KGS5YAJick3piV2qh29LBisFGUtD6yeyxQp0w8vmCzr6kGyBSP3O0SUnQGSnLT
6Q2tE5cAtKaX5zkA3BtnECLWAMl4zpjI0m8fNz49HwGesv8EjpX2Fim4WiClVOegHMmCau2Naq93
+nhTLzqBUu/egGV/ym49m3WCCFZXJMg2/ly4CW6bZ7uvWfRIcEhkpmfNU6Ic22a8DBMaiDLcrAMK
esJZrZLR4gzIfaK+Db1sTMqs2MNiejFAZ+qkEaSN05+Uq0eOku1VBPMogFizVEwsDQnu4dRGdcaG
aqjhIhHroMrtMx5Gj69NwGcS5y8Crz7iVege27qoLh4SRnwpB/8IuilTRwAfzMNqnG5BOhZJZ47y
1iaYnvj/9sLqQ698EYwueYLDpo4KQYxBxp9oA7ngOg4q96HxHy5oHTVTBq42jJe9MAYHxoE+FcpN
5BYbH2ObuuvOGR37NNeilfGRAVJinVuSZY60A7tyPoaDyFmRy+T1cc6O08a4BmjmhchoOM8PKSU8
p+0G23BAaEBDyjE0R/b+1RC3XoHQrrEUmip1svHM66PBHXXcyuiPJbbhqUFm6s6eocHm0syadHRO
fHtGrbJJkc5S28e9yaHk2BXdvOeVuK2m1VRbBsfQbnLGP7ceCItplAd64CyXr1aFsC0n0aPCuRwc
EaPY2eazZWB2U9OHpfkFGAdAPTT2+P7Hxgnul/uHubu+0AaZGs4k/oO+Q59z02xrFaNHOJuF26Uq
lARKkqmM5pv1y8s0vWioOk6Mr3y+2PkcAfODSNm9JDrQNz4opM4Tkyc0YfmES/WhB5nZa/biknuE
uMNcEmehY6vU4n8ennZZrbWXHrePjUSyYS+lIl+xX+joox3IfyuNVuwR4zVhOg3wAy0AbX9HgRRK
NdgOwB6H5dO1Nk/Y0hwtoRqWRnuyVjPQQx7sAkZ0ZFCPu21If9pdiwwXgokLQNdKNd/VmbE5b8wP
CGNpjaIkufkh0PRb9tTgmMkd5OFyqd1gl2bILvd8fyB1YtFBXbCMqgJJzJq9YCcY969viUisq394
MP0u/HGTCS+8adyPrtmau0vdP78XPzb0xFGsOwylPCga78ZotmdvA+Xlo+UQ+mFImNiaIdkMYJNE
wuKgxgqfY18lENgB42/kfB/aR4OVuPfx+qh5TGq1MrrwovARUmAqPvtz6eg/+6/RYda7Fg98gNu5
71TDDAwr155FOdEmqN13wtDq7PjdhrLF9QckogP/3HqX/5Q+4dVmBKXXI/fiIbahmsvcL7ZzmLUE
42AGQsR+IMErsHUp4BbYHUwfrhWiNVWU2InTXTIwoJ13JAsezfmcmWSVj+1wwHjCMoRA87g9ecSa
d8utHhlmg93e5+zm+bd4cXx0aNEJ3pVEmgj+dOSDYiyPSiMKZknBPwUgW4XZNkWqmgPqYY3fsZhM
qMgLen2RxSt4cKkJubDbSwWYQYDXC5uU8KGQUeScaeODRdmmL9ML87PH8P6rbNIwEfTps26Iiq6p
CvEz+HG+Saslf8V3phRX9Uqnphah9T7bFLJ3XrTHfl+hmpM7KWWKbmuVcnlXKFDCiLFVJ4lSIRHd
qWJMB+m4+YG6e3nwRx9oZWDlmyS10kfTOVIMVP3O6oiDRQjsEIe3bzUGYbAvEhMxcyNi2Ovm1t+C
6WgjGthX4SE4kxpA0ZFqLWE2KeNw21HCoI15xUDSzLJnvAXv3FduLYEA0CjI/QlP2oqhIajA13Ac
R4df+ZikhqzLqNNRjyCBQI2AK+hohsDRSB7X0acwPJchd+suJHHXs4TifJqVbKb6ksPAK0Rvdbpr
RAnc7Dp+T4Xh1WmGoPq5lmv0801EAguc/GdI1++T503MKDxBvLSVzRU4MajVe6tIxuV1dYIdluoc
AouquBuWiYm7eSRf3tuxokNB4tFjniBqnvgIfiS8UKt5caj3LqZiNg0lRY223NwUCHTMYmoO65eA
SmhF4MkUiVfh6BgMpotnHH7vPIXt5tCHLlbG4Kc8tr8UpbblFyfdWoY6wlO9oaFV501+FGt47O2F
sCJ+ybDHbzw/nZOZlQVtVKa6+72GNboZBxkk3K8s0SN2Jej/MPOfkpK92ux1azk0StNputJlyY6p
B6/QRLuXMKQcV+Y+hHeVvuXd/ExgrfTjKfvn+WRt15sLLfFCW0dQ1ZrTjqqmnjwdFaigXlnLV2+s
rPfGhe+zGbwsbUzKRJmSqxBOLFeNNa3UUHvzZDHdXzN9EvKsIQLjD2QvHuQqnOuTYbGWE3xbIgP6
KM4CkGf4C2/RQBAVnD3JnO7o4TOdKpPO/xHV/mzgS4d6jyyn9GYdbZaOeUW09KN9mUgQiMjrJuf9
cZREE++cDbITneaDuQSFXChQ5aWnIrk26ND882Tm+sGNB+B+93bnoa5uWe1tu1qeogExawUU+oei
70qP/Qp5FXKW/nqoCkhD/65mmPxA234nSwo9JKGjAgL27JaZGgmwnckMoTWH99D8aJTWxuIAroqW
bOKPiAnNr9GQLWNFDSIVpMGiN30LDUhTlD89Xm+m83as7FBZqKnFNJO5Z42OM6s5f+xxnp3RQ4Ou
EE02ATWUR1HvtMvbvioJF5qzT4YEFhmZv0+GzmQNTWw1tKbqqKdKcgFW8G2JXmuqx5tQQbtwboc7
e48qPB+9ieMEKwGCcBRUKagwdccIh5Gpu342uNqUVNlxOeQP4DEPpzvPep9F0DyTeqWtFT7v++QT
0ZxwJNOBCxIxG2CFbOQg7ulguQeypIHWikjwTi1RLgioG1amnVWoVBwRxBuWFHxaAriz1BaIPHmx
GF0Nejlef0tpoODgbbZD25k1H5EXDjXAXu0bFvMhTABuyZWFgAMtysf9lbTfM8/ZhdeNiC69Mnnb
xEbINiKsyjFdwzNjSLZvX+7b3xuCoJqxIOXSKT6foG/Z/pIb4DQvrbVUSjefsgh4ERW6FOpqyc2l
+L31dhSRykb4AMwAq3AitZ3gWkJt7/DN3t1puqsIRvGkAQJ+iS6ZVmjEJIg2+55jdiJmdCgKPQZk
oeVL0lrQeRQzwnJ6sl1XghiOhPMBRhCZCkA23YDx4brFo/8lVxWlgFuXH3s2HBqcM+qd7WZiaW4Q
rDNNpurwc6STGI+yO6/3+eGzc7qhaym0QCBIL3lqyuXY6QXhC1A/qxJNYeTb5r9rKi9nv0nZDHVd
0Q4UiAsm6fWZMpCM/U9HsDeGB9asi8PB43NKKizuUMZRsqXBwGMLuKaMsHe1IqjRbc62TgG9WH/R
jYtS5qKrJgKmmqARD86XKhSW4RSPKFpMdjF4BlD+SUL2K/OHCURGgpCXTqIq6D+q5VuLGZ2UPkYX
q0cdEd/3JgYfZH97F50FAiTXeKBJ8eLmBiasTlUeZk3WsxX1Rd4iMXage62QsEtN1T+2bjIkQMEr
mnYnjU79KmKWdDpHwhLeGxFriSzgycrikvav/TLT9TFoYKG0eNRWBBtWnmsAWBDMjDCE8hNYdHVQ
786R+6Ij6/67q8+SHj6VigZHjL+eGZLyTWiXnV1FIzitobItMEfOa3VGGDYRLXl4ZDCOPMJ3kNZU
CaP0JwjB+j8Gt2PviQmVomXoCWhS9e6dkKV5wzz0AxPZc7LWpfFQWxaIuQwgZcFlUKrbVdgb6tIi
JYspsBcBH5iMe2lfGOZ+8qPHqw9wU4k1lMLOggKeHBBn4/bPsBzHDwAJTG1alPL4rQZQzRokpnl4
tzmbTRpufdYzYs5/M1mAFhbTcVqtKSbHMwSjK65To4+MKYq5TodTvQfd1f1Vuaai9wafDajdeD64
mwInrsrg2Rz0uq7sKg1DMh805iO4BY4dbeVtgY1OPycQPH5MjD8fss/ueqEWh5zl4YR9JZ5EkbAc
iEl3gCXmi6mfz3oaantB1S3C1aEqbUE0wF7Lfqavi8E1M+km4ASfdisKZilWc1xmqgKbdTvKFsjL
r31glSpdPk59gOXkIIlaWCv5GP6vUunB1lCnaByJI3Sm5T3IpibYBuP2ILTjul6wB5Glx0U9Khbp
9naEMqe4VyGUy4J0j7luct1P5Ks0lRZnU4duDCkaRwqaAWmgYnOrHlAKlUv/sWDgjWjZrEhP//YP
30gGPyoNMxAu0Xr9X9j5OXWlRR5pFW6k2aKZUu+V+Ky34w0PISdQBsy6PmPifXrKs4NVGcDEZRH7
gk8r31emeM4uzt2BgO7lv7wBMtgcQSes1/4pgcim3zwoQUHNA0A+yVRi7e2DMmIAKYmExfCU6eXr
xw0PZap4kP6hoia34Bv5vLcf2bYzrbRcc5hmnaYCLx0Vhqq8SumDX77nwpDuF+eAsKJsAm+uHkkU
fElKUZpCXbXRKoo9yo4PdIOzCRWpwtAv9FbEWpL06fmMefJ3nsTRh8uwVIBJQJdPuHljtGrninyr
XOXv4FFWKZierOjTIUwDO4ww1JHRI+DVEuNZUEzrm9hauDygO9z4El4o3fwLAgqHWrtKowCilgLX
BwezzWz7UIn9Mdxqa0KMXkp16N2o++ZTMcgSSDuSPxfCErHsU5issJboFX07cAJGCRtY+uXO9MBQ
56COe8Dj1Tvtxt/dqfMnyYrBymqEP4uOE21FQQG9mqsBjIC9/mlvpyAWDsAJbMNZjhXuxb/PJJNG
Dcsoq5s9lMOyI1rqGaZK9UVxNIDKeOyuXYmrlxtZGb7W/F4fQGFemWrgTdXfEUxf/2HtSrpTz/VG
45ZxNLPeQGmQYsV21potovi2s7DtutCHCZothGxCz5AlTu4l49IcCPw881yh1yLgSU2pAqIr4vi8
o+fAejP4SrooxIHgkXeuC1FrcxYWJo3bMBq8AeKuhuy77HD3dB3ykLZ+ovA++36p+BCJX8WSqOK6
4LRsRwPtOCsZKH3CkOwgVvYbar2t2DhSPZL984Hte6fHX/Cqcc7cBBo1QADD6b/RAZjhncppLDXv
gDgSwjHR4rm5i0ue7rI+MXYwzDvOaxX9uYIaY917jXHVDCQD+5Q/qki0o1V8rEDIFQr8TF8xDrha
EPnzBvqRi3s29qdJDM3U+pVU8kBTpsxoMtrf0PmUniHK9lqAT3TcZwU6HQ+t46CrLY74JZkysRIT
aP2HbLt6WOmlhLAqu0lsCqbxIMtet1CMpj0SOqNwpPzaAGsza+U8eFk+dgvSuJe1uhL9p/M21IgG
3o0RkELE+HuANlIeka1u/BGQvFnUWAKA52aBurfSC9AzudFM7R1tA4/WSlZqWxHlgjDPczrslUZw
Jh03Yvy2QAd34truFtyWFR1e1lXvLltQQ5VnL3s1i8+kuyei8liNIUBc82UFJFl49mWx3FNCjw+h
0YZXvHGmae5bqtHnK2OhwmHimhFMzaWJgfyknIOJF2hjPEZkI8R51HS6zYAcgJPdnKzHfOpUaWVx
4CtQduALvzr/mcOi2y6v0s2KIaopyf2d9bHzl7oByTJB0xE3EhAqAWo9KDOKesW0Dwflb1HxddRp
EYfaUPG6T8PEreFXOUCvkSPrUJyfiIpWH9kXQOs0LG8KJ4reg4nLG6Jp9h9+S4XAIwuLXYea9+yf
Db+dAVqO0ZIGNySrHA/j++rjRGdlKRl1JaYxvvMAJzvKA35kYMEWNv6D3/or14NcCnQyvfTxJ/GB
ZyJk5FVHv5ZBulPfC430uG1r5PdAikwS+w6tHu0AgBU7gdAHjA7VirsSvAZe74yl/SF0ZE1VOJLF
/1zJFkE3BD225YOkz8JYjQCsc7U/NoVtUtLKPj8bcEMEM282qNGBZizKVRsH7cisTCeJw/nGzjiK
ZYKRY6Rut/ed0D6ClUxsDPnjuk1y1ErZab9qjV2JuDx27P30bg2cBPOOgzGzLrEAfRtBp7Ov9X7Q
KYHu1SpwUEz5yIaLzzWjEdYB8p+DN+LCyJVix0eoOJ9uV9UVyZEIWP7/SDrt2r5YAazSJQWWVJ1u
XBR3Vvzc2lo98XE+qM9jza+1hasXfIN1KCoe7OukaGkSjqreO+IW+nFzIkR4V+2RQF7uZfTMdpOH
IGuGlxOIY9mU1yAUoWP4m8rxtPFNKZWKhPGc8hz3kjGbNhtxZttrMpx+BXfN9QnMAfAcHuxMdWr6
uGvqndwydY9hvM0yDwmkXtMGOK+WtvZ4wFQRDLn5flgnYbggOFjvZwjO2zR1WE1MFGhbHYVe9cA/
OlfGVun/x/kqhcGCXf51nQ7l+H91/uFNfZ0geBxhSaRfxeuhS0524hy+DF5Re6fgl8VqP3RvfgIZ
8E6U+XqXfzF21MzEkBL6092hRbnSPMN74bgbX8gl6woLCQM7mCGUuXV9z1NopC7Sfm1gdQnXuHjv
seN0JpCAAKaMT0n2BUHOo2GCHjI6reH2lYj7bldKdO3catUMuYNJFQ6WdeLuU4cjs/TfxhN22yGX
diCvKO6a0zXQo1G4cDzgtvkRxQk+wkK1D3ecUjFf0FQKpcDkUL/CLnyeOC93PRtaOj0G+h/hg5GU
aHWLE37xO+hs49VLMHrJzSDVbncqRL4GwXPvLcQ6L3jDISkmjtHX+fsYRZw4W4b5Ju1oAUCK6kG1
zaA6zbDQQtqH44JNZCkDcx8jWWI/LeIOKZuE8YDjSUBdMSMi+bwbDiHl67fc9+Ur45hIufGPfORF
WtN5+lsSbQEFQSLLmS7PX4xpxe8Zpw6Nr4J7eLuMcNnt1iq6KtsDBtWeNZmtb9QyHjMHuWZiA5cl
ZGOivNtfngOFEzXK0VixWlp0iyI4hap/OnEil1NvlOBtekhNRD2OYoCTqcIm45NZo06lpdcebP0+
vD4xQUPWignR34YJGYcgvmP+GCXqQI7B2kb7jNSvjM4DcYBFJpO3D/80V9u87PK2QYxRK+No6MMl
Z/k2+JkTbd5Q2LqZlKX/aN3JQctg+73ZRgzfVRV3RF0VTZpsfuqtMStkzWh+uxMlw4v8IRlRB5jI
II/SHFsGpMED99T1IRJQV3i+csKsTO9J8MW4L84hnZQoZd0TlT7T36fuW/8R6JGQi/dc0+0YgepN
bZPe9zR4bYbS5kS8+slORT6mGhC0WrrjrYTFa/VKFrYMY5JSL9R6NrgYmu9IeNe17F4gkW10pIIH
jZNZjoHdOHe1k3i3UuqB1Y04BBYmcuqMEdkuQ7/ZNwqeLggdb3FC5AwdeokdB/0fFUzzAARzgauu
tml7mlMBN6YpYuiJ6li39FOd4JM4cWgQ3FeSwAlUcWXiw//JQnY4veomYKff4eeN4fbqMrV0xNlt
I95fd1ZV2+3d2juuSd7xYYO1BKaZWIvbtLV/yK0NlIWSV/jIrojkOJwOCgn9w789zC0mJM0lyCXG
wGMmNN0i1NNz83qSjJ6hKw4ZPFG6iMDNf0JhiDClWeeHjSF0m5rJiugcmend3ew8Ape3tkamfY53
5fiRIknXriYwL92pSqwZBT+4eGkRL2gnj7u+tdTnsOhoLQHEy1bN1+oh58/2HV2MkY1f0ImvAzbz
cLM7gJ1wa7S7UwepJF/D0GvnPyxMmfrnNFi6XO/ZP5M+rMWyEAWkJEMBieD4vEr+peDhyq7BZXwx
vLtXxrs9TindM0wMHAbmT5YA/ZHQQ7eulf1Iay7nXQBgi3yh+rl/e35qJG8WxPY7eFZbOvbDImBX
QRvSovFCKpjC2Yt0syEPy+IEV7JY7EFk1RWrXEx8hS/gWzoTgjCMX5W1OljFwotf4qT0xRkKSya4
mP92d/bi28wZixsAPCCogNL/zpQtUWNphSgmT+D+2IVj3AkhJ7nh7jaYGfv0FKihbrGrwPig9K2O
o2VfhfY60KMpWn3e4CIJnuGZ4R15OOCyLO2O1GaZceTU6D5d1/PPml3l/uOfxK0EVtifl+Z2DCnB
h8gMhhM8qeL68g+6Tpnkeggr8W+RE3W9ZKDsemqIQdFp7FRkVfCmB9BOSQI7NagGLeJUylMJixyl
70K+xbBIvrMYdh6VyQujyjA1UZh8fBHIkSEac1QCV6+ilFYQahiC9rmrqxPW3LQrWhVt3dL00+b7
hfTOO2zkjMLRr3CEE4FhErxVOQqv9laTc1P3rA7UMedIIJQcmGs5q4NZo19Lg8Q5kSE28DmCqfvV
xrKGwwYOamG657sbnhZjaf3aAxa/u2J24LhUjt9kHkUktgficEwHnifwXdn7JSEdOW7qA9vM5B4u
IuFYZtdbppxXv8rjw50yiE9e5lW1H/99YXUbmPResc93QXS1QoDcdAhypGjHFMry6iHkndbu8ET1
sa46SgQOzHpH4XQiXLRfq417gk6g+EmAqzpzKp7427smp2PuAlCVOWI7z3K0JhBmaaC2stN+O7W6
6Rhi4pWbq1mxJRCKtlJ+c7O60XdJAsqM907vZ3AXIHiVYzTXqJFeGWrWlgPK6Nxc+jVdd8CqG9/0
EgBvnrSa0q52B4TeBDT5/uymOfHdfsE1elCVndx3DgG7ylVuZQC3OzYQazvziqTPHtpaonzj9iXo
CW9gnXT4gFV4Ln8NFnofJovwUQWUqy5X+PfhsK1C7HelRNBa3UsTBQvNNoAX0cUnYsXL2E1ShkqP
TH0hyxjj/VhTVKEfD0kHie3Wzv3hlIVufDT2D8NWCABJdaWYWWVVkbCghYsxhL3R2bwQ2HrD1kCE
TF5WxsiXA4SLG1tGB5oHL0CL4f412GP1jNEItCU3+yQrQovdPQP0N2U2tmp9G4Qsj5BVzfZMM2Z0
y0Ac/rLpLAUPr6rzEmwTExX3tl70U38o/H7YEDZAcB8bKJ5i8KXXICQFSAFgHVPp2beM5zKT3B27
WXRvxE0Ix+ylT0crM1ccUcQy1WtAySxn1vZEje8AHBZaNK8Ck74+BE4uMcmUlJUf9FjHtebJiBFh
THJDPfoOTS4jB2Fo80R08hiHzqT4rQ/vTihGfzQr7URmpEbqa3IWiJ7jFGY5V8SUWv962fexhnIu
aCse/hL9WYMkFto5zTaxVaZzhs6GgnbDUFS7EMuAafvuqArwHMSLiXKW34Gp2Fd6UVEWYNkLoza/
0g9Iamcy7Mipv3+kgWs8Jxn35juxzRK88yhaUq1rWeeLF9QyURzum/J8NE06/NRYYiuxfBYG5748
MpObiWiHJzjdgpfkZ5OZFpfoJ2f64IkYt+HL/OkrAhNF5Wl+mKGdGyg3OeGEC+m86DwKngOTH8Kx
1UyadyCwZYd/8s+htd/B02kbikgNZ4MOZanBgLRDe8eFSY//tIfCWe+L6iHJpeqXXGNUrOvMVOZb
ByKXO81Gj2jvVNWyu7fdHaNcgNHpGZ7LtsBAbr+f///ncRb22MLeYGgrXJQ0e9quEy304+gNZmRO
WglUGDW3HHlv78BSWPAJiOS93P9hdIja46KKPgAn0RE07u+J4UJJeMieBziq9DfLKrUZba7ICJMT
kM5OxjgukY0JPAkDgIs7Tc1tRvO9qWR5fkxD40x+hcWPGQoYPqCRq1/qwk3+V7Z1nSUY4kquYvKz
G2Jp5FCph/S8Sw7b82ka1k/cRrz3y2wdN2mLIqJ7QmR6hw43gy8sKKpQulhMXWWDjYNkBB7h4B5k
aHcTjRuklrZSJvIei33K5AhaYfICuF1i7oN3v5LCAj/Wkrkv18TpjVZLM9uEk030Zi2hJkr3BjNf
GVwgk2XTcuIrMqb84F64iRSvWWPHXND4JQs6CU0z2csqY1r8VtGKD862kxqc1j7SLKURK7jHaoDL
c2c3XlNd11KttluinuV8+PsfyVPeFYhJO7pFWPjatRdbDyjiVlPkr+H9ufwUMfpIHS/fQICJMHwN
6HvZy3dSVwD6Bb7hWCPO25ayph/yGZWSa3lIv76BNcoDSPM8rnxcDIjrwJ6aIo9QdfKVMzxNmyLK
luxrpZmULMuVJRqPYTc3GDR2ovz7eRMp8lgBZ8bpN48ykGocRSlZQvQin6GAKjZghF9uzASCtmKM
jqOD4Va3s4rMdagvc7TVXnjTiua4s0MIKpw2cbAsujCIvR/rlnYr4V2WKvz9fIOHZhaNeu2uFCsy
VmdMIlTiHKWBPsEjc3Pb32SkJh5kBCueHQvHQdk+PGZ3j8t4bFw/jlIWIhhWAVEnP0WVBs/Ydbxw
jcVtnti8Kaa/QUiZfVZzZQsoKAXco81+kHbX5/HQill+fKbccNVM9X/jKIbgpLOcGpLyQMewXBMB
mVwL43yMoIQNhM8f3TM9EyBVPuiUk1DlLqLQtoJJ/tSYkpHZif2hYg2d7FozDp1XZosRO4VjiniB
jTuuunxLHgixFSRXrH+9s4aVJUHFDwAMRcEb11U0sIss3yi6WJwOvTqoejmkfnyoPzUWEVCRyfIm
bhuGSDLphxnu4vTAfdtQaarkawesPB7myWTqFSbSsYPqEKp0f/Ohou0p9uYvMkiJh2+77pO0OI4p
BbRNqhMqqGwCdS49F+DBgqBjZrdk0S5ZfRetGXTgNopLg7dV5Ea9KCW2dq14UiJl85zzNqt70LF1
kuzGbSzKBxkmNoVYN+obSLvCGlMmmdbh7SwH4wOTyluAAUsJ2hxpXwc2o2n+Dj/3fZNP6+shcDDi
XE9aFQTg0cU2M5xlV66+tDXPBg6EsKxQt2b64mzrytsUCiVNNPfBgmwTQDt2vMwy7b3Zd3XdUWyu
Mvxt1+HBRh9TOO9RPVp3lffl5Y1lAitaZNQToRAztFdPNeXF/jH0FKE/U0N/KFvnEPv9KGVG7/S6
wmHXmuCv57PUliNymt3oeObzVCgn/77oSOtD61VjM6EG9/SJN1D1eC3Jne0GVhtFZsyeYNpM5Ax5
VGXLhRI8WOqrooc1DkRiq8cNd/595D0fN+1DHzxp69tw/7abO20Q9kI83jLPNL46lzXVnY9geu4W
1XN+JPe/J/ywI9MJQhdZ6UmFx1k8n4SgEVeLz0z6uA+h4Fj7dD6zw7JgBXhyob4A1FzmWzikC1fg
bbDVsfxk+2de7v+6C87ZroVpj/seGwaXnR0lAaQI9os7wviXfUUT7ilgowdB6aeuK+xEO4NiHFOD
hLybuUjJwrtAa51l/L7HJmcmCLjKZZwnKj1tegI/7BSGmYNVpTRBmF7nfDpi7mPdPTAez4AzH8jw
nF99DeKZ3453VFGP+ryp01elQ0G2WKcUKBa74nMR67CSTdiv3284cX+JCAswGI73n35KNj9iF8uK
GrU5UA+BQQ2ZKypNBcIi73U3t0I+W/5SifuHcEzbPNwBuO0oqWIZ6kNG1ZpOO7lZ67HGtPaB1LmY
c5L4XFguOyHqujqAA1dZdNMImsYvIJ39mDlvW14CppdsaaehAegkcs9jecgdtYlc1xYEcsMBt/2/
SQU1cIU1srZOrR/eLgeFqDzm9fmzZQE524dH4umix/+1431aMYDyrR//KGAlHPe5EcYq/beYpsZj
PQi2I6XNuiWCitWPcib+VFKWGYLm/1kM+xB46F4pch2lZKTlFeRFa9H46r3R0IGsTqe/BKO5PyCI
4y4+bdl2ZAdBafQPVbltxOfHz+2eOJoJ4T2kafKl6KwkDH9s/JZxFBgIk4udY5g6JXFKtNbiZLnB
eu9DSpF1yB6MM2OtWRaWRCRDSf+I+HI1UqDYH1nsnaCLqBvsC6FOJf3bvkBAdewLbIYUiXaVAS0z
dS9tx7Wh1yFFKAGFWfhK+LyHs+CWLh8ZWEgR1cc1xYFMKzgKz3r+1dI483rTx3PgOqvWGeYf0b+e
QcYIzC/OX5QdDnlXW0u7tF/i86zXkknPmq2cF1kfF064mCyWX2hc+sx83Yl/cxKmLBJ3vhGSZscX
v7PBVdu8h/KzVrjz5FhJ3E9p2/MUBdFU9MjugjGaO4KhARFBcCfJALLjbT1opjzBuBgJPqaGkd/a
HLYRkqWjjFonn+txchcArtEIDmx5v6GmAhYBYTTOSkXpoBqZ+ZmQpuR0bihs84z8s4MtPR/+YG9X
UeS8gGhnCnpPY/zQN7ekMnOPJkuYECkL8fhKD2idU/EAY0o2aqx25sTSn+saj7Gc7tBj71PJ8Cho
MgngN29OJ7IjmCSzPQw8Ao8cN6Ia9WZCtv2yzwlbYCDYUmknJt0ADmTgHYxdrQ9BzTBxkKot/uCG
c0gNCG8Hj6dGYv2o+x6wuDD7uZ9d+mWIshstHo0R68RzV5n6CZNEVlUM+xEzGBzl7xVX7yoyPZM8
vpKdW7hAToz0od8YD0M073mCD++5inSZZo2wXb+fnlljZtung31/5FTk3aPEZ4d3E+JYCdQIzAyN
3Mcf+Vp6TYfYonmXSTRarkmhpcDCK8GOqShEe7eHsot+vvimuVoT8bczzSzh1WV5imQmBV2jMSuW
w3jbrOIbwqX43CSiuVF8sbimkaqlF6HpTSVNJLvsbWc38tbE9JIam3Eg4fjKyvrl4tOJvIeCc3lu
zmNaujPovJTJfWx2tKSMUDfxLbdiCSLoACAVQqmZUhlHdPkpHHB2InNPIPZHDB5vcm23h232UOG2
ig1WiaA1BchQXamZcK9A+Dq0otcWSQzeTKKV5tU+FA69kLPRwfHdH4HApLm6tZ6jjJs/WBMs1GjJ
/Hwur5j0uNH4iSlsLcbYXrFz4AqQZMnJhW1oO3qGOXsZYsIZ5VGdcwccH/cM8GwvtkXg1te+SOw8
j/6Lf8jb5Qbk4gUZi6sjC1TDivUHp8p+cxdW+5wSzWuQxVPBSgM3MM/A1ALh4ARkl9Narqvw4lsy
c2yS52PAjaWZVKyarNMD/A2fvXizsG6mba7bPSmG+RZZ9uzvJjBNzRCwtMrvy02cqDbtp/MXyTwr
QNpSQ8iJNJOgtjzf5WpiHCBpB7dHTd7vRvdsAHwh4wKYHu8EJjKs9IY/T26JgwhZixC2fd3AM9yP
xw3k0UALqOxlvxpDJ5/dPFJZ/NVY++D6L9kknUPrMOQJpRx0IC6xjFTXmqG0SqbWOObvWz0klJVi
XBXp7o5DYG7pA715Y+0vot8IFHU5lsfVCXnpZHo6QAKR9bA9hHE8qSOb2ZZ9ciJM+/QD5SGD4MJe
7r9B+rhr3BN0WzBPFljzHrTzplGaXXh8VaN6iOCKoySNLcez+HatrT8MFegSeLIHhoNvv+XvG+4S
TWthTZgl5LWdiW7sqIfqZDf86dhXB5034N9ldthhAbl0q6E0c+LqeV2/+WQ2Md4YVS4vo0vIdv+0
wDWzxuZzeCYay2lbAuMFh+XjF3ZRzV6zqXkRG43Vf2arWZQ1mBa0zuOCiO4qS6FnF2pyThznDXfG
EeooB7axijovH0EkJ35ZhdZE2rdD0XjdOVpTaMq/uNx9gngkhIeKpSOFYfRkf0K9SbWwbK/dznFH
+T+UsplwJUwXhOTpysOHMrh1LGkqTUvR8e/x6ZlxEAnnWE8687Txo8rm3ZROUN4MiVH9BiYLLn6Y
eKe2cPFNjE+FbdHx/3Ri6DWFIoNwojGPzyRiqt0T/QBW4nRuafRelfuzOnKHugyjpe8Y5X+Jr4FN
ArYEz1VOb5R2qj33ThlbkVaCB9bkXw32WrFLTvGlKShOfrjr4VoVRC8TksfUMUbpQNV3rQpvdJ8z
4LTfQfnsGQ6HvdaDGj35a5oQ/86tmnCJdiCBjbtiUoXqh467iOs2Ll5MrXk14hCSHcPBrpsOXbaX
o93gpFlvOCZwTTucPpybnXjdlCXsX4FsIo30eKXUGTzmmcTiJuC1D6uQRurRQ0WIx6xQ3sF7wJNd
dwVbn+mvV/tOQrXLyEY8DnP9GWtdNatTX5VeXI+aUlzS0tWXe+WNwY/5pUCrni5mnyp0aVLYSq1+
RbmTA8mfddCUsAMw5gK1mXnoKYbUI3k/HMC0IAOYav6+Td6z+GROVWHwcFB9Zdrycs+kIyNq+hrm
FgOihZrpqm7QxopRSMl0XTHEEPPYly9RNqZSdVxZYarXJ+i8ajzjKg4TlbLv8E/DcOJkUpAt36eu
bubbWGiE90NTExgqszlkXnaae1fvtt81fQHEnqEJE3/cjeA9y1XR0z1Yuw5sw/5HWna/+ZZ3JHUF
KXFCZhwAh+GneubjeECi5nZcJnwKL2HVf7iMPVeF0PrEbg3H79pb3hkiYLc/CXrQpvZniddV/u2Z
kTpQEYz5rAMAioRiDmb1upi7KUFQmWqsT3fc3z9e1CX11w5R3aMIEoghAIjil9LFrASxvdUWnSbH
7Ykyk2UAREBSz5X6tp3A3SoLgRSCaprKMlRCGsDFNIAxOUfxMc0HdzHJdwrIsjgfvFq62xYMQqPL
XjzmOkc8VBvlhfipxN+/e2rSCSZmQGOCwxGe9xXghn2pS5y2OooEK/Oi3LGgRKaV0OzdhyXy2piH
TaCuUjiCuWtXWtw0SHRtfagxcwk8pjwrX91keTI75McVWRf9yYUhzuehDeslTv9Fn57U5RkMIpkP
lelNxitXc9khU8dsTRBTBWzgfTGasePX5JbQbiHpmILUZAZ9lJcSKNsyBo8E7y6jmr+aOeWO7RYx
SyjTaKaFEfQjjUA9/weATn3TebYae5HFRWWe7wn+OVbL96lXsxXawIjQHOE3eZMjnasCnaK5QMoj
7Ch/ksAd0p9ai4WLSiYLqbZXsUWF/TK/Oq4oGhdhgOdf1q5dhAJPnoAVI+cx90N55GvyxsNnPRXg
3YxW+LnnYE7BYWZnmLvBFDYucoShTERIy+oXANxZJPCV3O9nFnBdcvZsNvEM9VVuSeIllAVGrfVq
iIylj18b4581Yt7AO3nz+RUP+xeHnetpvUKopr0hjMK2ofCgzOGa9qrvTXfkTlhAa2z27IISAjzJ
qLeG4sq01q0ZcbO8yDewFLeSeYK0NcQgdG9qMRgm71YHDGw+qv/Uwk547+zfXlLzvkroMRdQCgTc
+acSwXvI9bq7OGxGl63mtNpWuz1wHHU4QT1rF0RP9+iB8VifrfhNI58nyy3ssyeJKdntsxQ8wT9B
0EZ8PK5TW7ZNaFq/Rvqr5uIBbpRSlIgeti8h8qM+dMficxcA+BExrlzOsijD2bAFwR/hLxFrsHj+
lcAwwqeLsLwQ6WAeGYzHRIY8bUUKKZz3NRlnq5QkJitRjJAaZEGNiAuAZdhsy6+yNc9LqRoCklsU
+n0gU9eNiDDFNA5MOKuyDlay2807K/rVRVO3yvfqlP1bokSxXzhj9a/52usxh6yUsOlSVkbt+Xtc
fp5CDfqINkMCycnzGfxrn459e69WvnZg8jcg9vQM14SfPS6JDPTie2H3/MT++We/nTRWtim+4Ucj
gu+Bt+2dBFBXXyeoORs7Q3YOlKrEq58spcy51/DUE4b8YoiZCrWqAXJNd8NqZzRb38QygoUVFZQt
91guYLP8QWphIkAg41Ofw8QHq4okGvnL1QFhWMB+ADtsg9Ggteuxi37gPtR8jRAAV2xGPd+nDX2y
fPmoa5nr5kD4C1Kk4F7G9tye7qXT1mSe14+7SJ7kau2pfZNvv6GeXFm7cDqngWDoj8yOv6ThM8Ud
p7JqOXw8kD2I5uxBZGrTRLxLat44vAiKxkYUutV5pDPXdtzFUE5hKq5rJILD4dCelpqjOEhJhnPf
HksytKwmHiG4qLqQw+FpHJMRQRfQ1sVF39MLdH8IJg8GNrAGDtjzagX1hDlz2Kp555DV+AgSq79H
A2W9NRlrB9oR6tWWMQQytDHCBlwUMyQKJFopuDTh6ugVAslC5tLZu6SKg2+HKPtmDnOYq8vyLRzL
XIKbboHl2J2W1r6Tuie8BW9ChjlW6LTrfRbgUkPoPWpJsCj8Ouoq9rcsd4IQgcnOAzjZEZf76Zpx
wek+mArGmyaaPnjgQ34hO3XWDd0Mx1x8quKtUJatXqkpa44FssbPHAblOYgL3tqJhj7FFi5cF8Fv
Bsm7wNxz33W39HPbX4mkY1WD6R2l+fpTnNOjYO6aYPElWBiUp4ZRFWODDW0LH5SY+iEr/rF4TcTs
JWBKpXH7dHxCFRvwj+/GcNEj/5h2YkiyfS27glBYoUmxTsfW7GlqgrWlebKN71wwqLKkqJ79HJkC
/Y16A4eMHopsRzbdGdYICqGPh22CfaXq9L7EHmQS/WAIPwp+w2cCNSQMrDXg89UPddDOgHONbKn+
PqlUGVB23ssjAAvhDCveDOQafHhs4jDWsCFmgpiVJQj0y5jddWVwar+PlDJKbJhrWdDoCLdE+RaQ
Bkhfk8sAGT7Iqn8TIExNlcbX+E897F8f1kfJ9i5xVrbUxv/UT7078As1klFRCGWZPf0GagnrqoO1
v4tNVcPTdOnO0ppT1lQLrCQSs8ImwYixeev+1x992YqvngctKIj2AHvUF2Keq56A93tueBsvnjD6
Zzsb+r3qlZz2MPAt0DMBBfKRn+V8r/qOhPJ2IuwpF9c6m00dy+eW9sGMQMgwb0vb1dEQb5sNlxu9
0rS5ZTJ3mAEH2el5ARfFv65B3IyviMI6eqb0CkHR9W5H6k+2zAKXMiKrnHd25UnVBr0HJ8V/aQO4
dnxiVWXQ1Wi4O1u44FEurSZCzA7CN3O7y1E91PI3G3cvx6ZMwHwryvb+p7uMjAWn1vHu7J5Qt18o
B6evlE5vzfAEBVUhLrypnPzn5d5VCR00597Is/5RkYHbo06Ap0Df5mB9E0AhLXYzWM/1Cb8i6jgL
5tK5JKbjBSp9PigFZe4Htl+L0wuN3OuMSUYvmL9sUGkOjS70cWpkhItg6soqTATy+7CZDMGCiI8m
z96zvv2CGCudaG7kWCiedn/wqTpCixvjaklkBnM/JI8gXUM5gLYX0Ohw3Z0VHagIak2iFXjoyr1o
HGS75D+zuSO4U6C+45mb1cjJMPp/O4AxuS1Vw/RRHRgMDw1Ohm5oBukAzMXsOqvA6rPPupUndZz/
0pWw2EzhYDwJf4kDPvOUFJBJHkzbnsu0TKcJCWSskzFHg2GVs/4py/ZVGDpu4Wt9DFZ92hilW16w
8j/z56ziQiwZkZYWPT0R2x5BdcK+IbbjONOSaABm4UL188gJrlQaUZDB5XH4QNXzVUf5ii+qbtvS
c7W9dUeDSk41wSYFxWy5NEB6+jinCgOATCYfkSQeB6y7jPH06917+GoUhdn4GHyjg+hCkkB1oHIG
qnDIsoFzah7oSTrY8GLsJf4YDwcU+7lB00IhSNcJrPYJknBubAnorRQ2NLcz/pOLIfLVwjnDU1VO
JcmkgTl0Tm356OfZdaS53i0/JPGBtjyzaZK1ARKCXKtpuE9dT+xjHdp61EGGQBPgnMw6JG5+Dpny
5Cy3MPIpujI+jetAlQIIrO/HJitezSPc+kL4UvQgkko/t6YHXFAAAEup2A2vpqzq+RlL+kIOuYex
rE/ek011yG12r+Gj0aDQILn9Tapf1GBTr6iuXPHwA7lWJJoIOh9Z7W2JmVonJ4/4QebSinduAdSg
3/dEHbhJqxynU4bJMqLQXTAI6KJOYzSmdfXdFsNT1kkxx0HrAoqzckCIKjjvBwR+xbq72qLY30Dn
DqwzU44e25dPyRS4oFnNJ4t+1f0NZAfKKmDKYKHw07IJa7RFzC582aQ4jvb9j5z+/AMIUJScsXd5
VB1iwkP8/PfiuXli3DBN9cJSYmCOq1I5ZvpeJlXOhaBz5Xr84yAM29t8jprxoGnRX8Fx/H9vbTQh
7Uut0GGOB+M8Q+gkem552/1CnHlawve6QTOCWVM5V15J2DrOyACSt2GGG16Qk1XJPnnBkjjhx39G
OCaLrzFWGS5y3o235lR7xkjyzzngMGPhyjxtMsjlxv18ykbe799Bccn+kxsAzSY8QFKTzVEY1/A6
0G4+E+Zvx+KbMANIwEOh14Vg13CSMEfA64YInYiR/C5MeUnGD/QMhA/Rk+W5PL6RdeTFMkDYjoPj
dwmedkPAg7CQcXlmKRFJpGaI9reGLCeFxMJvdE8HQ2oNKZQkDMIIHXNFfloTJr2QY7ug7/oZhdMG
KpykDEFCDiTX6kYXQ5wKCIER60o/CBUiHrCYOB5OakLUd6SyCVB6eN2qL5lPRx6URJ4A/wr8cC6K
rj5CDTIeQY2UQP3LqHcWeD3x58PtdGXEB5EYNOLyASowpjdut9YvrBzRlabZCUlxzJIk8yVC2RZP
rJt+jfNP3zvU5BUB+M3yccFuBeKDeEncg87hCWUGV7m0JjS+DxjZ9CFuOHBhs31uElCAYr1LMITO
bvQPvn45VdziLBgIrajISTia1+eO95ISZUVsNiiHZhK0e5HuoEmErlULq4fNkNIzM7f9yR7JDp/o
pU4tbLI9IJMByivtvgn//sB0kMYcHBJYJ+xVxrLDJjReXO7hFIKGqGhSr2d2vJSYllhsouPs2nNZ
4HvhbDXrXtz4RZZFXn+ZPGLwqa1NbPYinJTCPDs6SN+aKvkZfXOxENHMUIi35Yoo74j4pcMyl/w9
rzXO7osJk8VrODlWEn5UQwlH+wB6OwwNUw==
`pragma protect end_protected

