`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
oxTl2+fwky53hiXp9UAfqnrchlduRNvzVAXaNi6sWYQSMfmVo3RXJwc/jpgk0W3858Tq1oQkh0xg
ksAtKElH7a83Rb7lBJ/mhKHi6wXm5GwRNT+rgbkWj/TOcx0emRq9c0wSf4uU1EjzW8xxzbGyXDyK
3cfxRGxcNAJkq/WlLsgzmTGvoqxLADTQEm+qna02RHEnKBWDuOIrkX7MZqovr0oBge9U7lF+I2o2
DhDEF2O1N/Pent9AdPBGifvI1bcCiNyyD2EXtdOu+zfgnFvp3meRzL6X/XYrJnqAgkic8n+txi1K
uJAnc3SHck98heWz6Rxv7/JzkPIkAp0Zh/A2bg==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
NypiSBDCrtZs63g3i7BbRzD/2k10QO88V01yezZuuSqEOnCq+mcYHJpKLUK1FX5vutZwVn7ACjfE
wxgF/J6B/jLoXgUAeEvcj63faGAPrX89T4exvcxIqc3W7wjd1LHUUddoC7IPvQHVIGEnIMqKkMpK
q1wOjjfJrBQIBfwJ2f77Pibxmc2TyafKf8zD86WRqnA2Mdi+SR53djiCdKR7vNVp8ORMWc5Wdu4z
l/f07hQ03gQmBNk20QDw54B5AN5b7K3ycYvyDdoE4tg56y4MZySCYptMvui6yF7sh92Q+vjKP6Sl
FvYhEpkcz9+zym5dkw2Wt3Oer85N2+uBScqiFQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
JN1eyGpZfqySkRDDUJo6OV4xMRbCdGTpy702Xs7eBRFsdBK6olVsrY5v+CQmmkHCTNO59atSgMF/
fCTFjz0oEg==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mTnwPBBthhH3g04Y4SBttjyj30RfjIBtHfp6FVmGM7w7MPqYu49F28Vh52YEpgsv3Mcvl6rZVmeH
vOcNTmnb7674BAgZbCMGnsQ5LSrgq/QFGCQJvEo2aFrClxP50dcKVKjanmhGcJBlPP2sbnj6sH8+
MtjNtOWv1IHrhxknzSvE3cmn7nnCwKku0fFRR5s8d2ht7lnuuPTI4IbwZx88qt5KRhlOyZ8ypmHy
ygw44CQqmYPhb7UTRa/+mliqZ8XSVIvrldZ+UlU/mriwltviDF0BJa/GHo+E10iMpe3Dlt4yoaR2
m/tuVVWFsI15zjj4ZbuWRkXHqIFBlsa4lQASaw==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
BmLUrCxXQn+QR9d0bwY9iQ2+yAVv2QEHjlQfe4A/gnfxPg1BEyIonjouFFiCnklBNK2ZQ8L0CWQn
pC+7SQhqqx3kUMIgD/yPi8fBYzfrQ9nFwp9jYdhzm3+DqOaI1+iyB9ruFbHEvSGaTK7Qk1bPRmal
w8iSTXjer16tiD+NYVtyJ5bPBwQi48yRD6By1jK8Xspr1KuDs5cNg5LpUNiMkZ0EmH57EyC8rCH5
PzHp86LyCfs24Li3j+63hnXPCB8IMXbRe1pyNuC+xDI8Erlh5oW7eCNWs7V0I62SyEM9Dq86Q3/f
y4h5jHp9l3+B7mcwckI3ViocMsKoZC93h/1P8w==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
qLALCB3FEpS30WFaKBXMhBX8KZ9VGFPamJuxJ8GUtfwvJrloxrRjzx2guH3xRISmNeBbySD3l1oh
m/ADuH1L8f/z8Af63Mxt9F2FPXXRVFBfPKEHAjBsXT6JmBknbZypaPKTdLUsLT8EwPM7F3C5AxLj
F6C16X1hUmA0InWRWjE=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
DRW8Y29KjP5L/O+w+bxRIG6nymkrMBlaFZ8my41wFOhHTgD9wnvUCg0y6/kpLsKAtoJSsEfVs34g
HxdvOKc+LFDJeFG4VUpD/rY7Jj1SLCS/yf41qyE72NY4H2RBbGenGIAQwsmUkwuBYTWkv/p1B0rh
8mjqhU0PSXVg4Y47NUieVQjKxfKFx3ur7BqhPaBjqysvVC+iwJhMDpEv95KF6IK9ytfGfB/6cAGi
HPAYx6vT2KJDvrmCflEHms8z2aK+4acr4Fnme10sjsXHJsfn2/i+WMyxcLxaz/9kig/ZUx4Iif4A
A7NpkXfqerA0A+XVGT0oq/Z/pnTA8aiQld8Tuw==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
24JJN8iMi7zuy4+fOsZPrTx2I5E7mMmacvxcWIp39OR3g2or4JWHBbmfrZr14pCQ0M1dHkCIeW+m
bn7fW/Ng5otJPEhVCoroKct+4Ey/vFB1o6yXh+bjVRo7rXoEqCKQ9K6GXiGZjZBcYjEP2Am0x9da
z7HPepMoUMB8TuQgrmYSeJWBmXwJxkBkBRlqVOYkwBFfU1CLW7aCkeQa/XuIhLHHivp4O69CtIdC
4/ukZcgs2UU8kWbF+TeTw3+z+IFcYLw/d4QEr9jkRkIYqmsEJ3Duc4/FHVZI8IG8cMGAbq4kd3s0
knze9sPw5sCg8dJxFGEUkw/iJzqIPAtj8fzcuQ==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
pJXC1i+2EK2zXaXJvvTZv7E3/f8P7SzzNxhA58aOu3SOWJYabFD5GsltMD8a4SLIDfXnJd4M/+XN
wMHBxpvvBVtFulpvcvLeHv56zj6PaF4IGXLTZLsLDQUasYCCJ9NOmsR8rzGY74vRvVqlJYziJKFa
mCIURKorq3qd1Y0OCaw=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
go6N40vWEFzcw0FqJ12M0F+JHCjteoN2C6R9cr/ckczhelRQ0K+rg7gJAhuukPmowzZ6jvrihFki
0CpCXkN9o9/kQWn0p/2RbrPyICsGXmcP6epe17zV+0d6qXglQQbnYinkacAINXtyOX74ZUTukqPf
cWcFoWPvopRpzltS1ZlllsblJDaMVDdkffNN4yqj/ifw4JGQXllCxnkf6fpRyCXfSy9q8bWgcCsf
jd8kDkHzAkDNrKY7mdiOfvCFKkPtUx9FjbGeM4lmrNCfMqKOsT5X1PuHCiirn05WAh8SpwIGl/AR
amVxRmKVHOX8YhypGJ+53KaH6cbYmT7NhApTzg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15632)
`pragma protect data_block
H0lhcNyawur47m+CBm2Zf9K2aU6RgL97WPj9q81/mAA7MFQ9/QMYFueXLYSf4LDCHL/JSwEyrqWo
2p4IJfngQh45r5ySoMObEbZxqtSLi8kLUxLgD60wTUdaZrEJp2ngxTaJDxNpxJ2wmDLUhlnkFe9k
zEvAuUxmJmT97GzUN+DNKeVmPASQG6RmN8nZw0AUZ+lcI2x24O0ZvWBew4tFUuJR/d7cl4hr9dKl
NyCmfIoTW/hPpSLPWgCujxfhLM7tiTvPJNc193tFWy1SFw3zHPLC1HFpjCVeqjz15R96lqAuaan7
Jqu6zlNzxZ4cXq74n8MorgY/9MMJBmN1NrSvOlWQyoU0EQmo6lsv1sySjoFuWbcuihsqeSwI9sdx
YFqUhMHVA5XVssOaFzcBqrSF3J9f4zeRIa9VtOR95q8b3LL6kVw0YOIsXKGC+zKZ2zLPOR8lBboQ
oA7ziHWfCQxdsGjxMmcvswFea1uGJwoOaASvFkzWEX8A3Ib7LBo7sFxkH4QVDcFxL3ldE+IhrtM3
OQ8CJ/rS8ADQcyOGtjCmGWzQZUMdzmyN4TIpPCAS1+ld8xBBqBANYhXkKbtoYJCN4FH/qI2ayAqN
sKhIN3M40PvGN5p7Vas5IC9/WS47yKJJN3Ok32wYS9Fsj2GogHAErPD+YlXKp9rS1/Z0RHpBX4eh
7rPBuUXIQ9cX+ARPzo9ymNInhPDHcRfAMJUwICKH6TPEbqjtz8cXybSL+ad7RgXJObf1ER4gUBJR
eNS+hAQ1VaL7R06y+aj0DTyaz9NWdMtseaKGtLZKsxdrIQYSaNP2uCrgaPoCZaYN5J3hWCxZr8Y5
kum5DIJ5OEV5I1zrzz5j2NsaNj6mERJurn7DlOy8UKRwTbCIi8Q+ASrdKJosyD2HAANprumsHBBT
GWKTosvS6JJue4WwBOBeVd7ZQzZWbVUYSePlbE0GGnpn2Mg+Lv4HJQSVIamx2AjrEeBUZEvs/vYb
3aehF0TbqUjXtwjW8I+vz+taH5MfU7bWksrIXC/G0PYCN6RCrKWh4OhiDH3uURIopvwpPVnM0QTo
66ka3BuyvUOeRPjQvpqDp3zTwhMR7UuTyHpbf8PV2t8y94k6TZ5KugiGFcNa38AGyhQL6jmnb8ec
cPt3eN6Pn3RwoSv253wGevP59XkOroCflYyDHCompz2PDS0cZapUQd5YjRAF6JfN04nJmqCw2zso
zhJCuPx02GNeesxBJ9oQPu4sZOo3gvR9dbfd5v/B76wzZu9usDDfUOipKVTuSGxWU9nq3dOh3Qfx
MiPy6ckmDbrfmgyYwLcN35cQzBSGWTcCJeAJoYcGzLWCTEKWSr+17mn/UgGmtOUhT1B7PPv54BbY
tirkcnxtuPwhlpr24n0mAR7b3y+NTCl/Kv8ln4rxzAdqqX66lV+oN9k0nTg3f7soSpUvpSLkUCTQ
W3BNCQB1RmQrsuh82BCp83S/R5/a5/12yWRgaeCKrmuGxnb202m573mfKzPlAKvVlv5V6hxcVwVE
w6HEWQ7zZBZaO+mJCfXdsjd5FfrqglOsnzIJM1nxFARL2Jx3wSnij2TfCzukyEZN4rQviDq+q6kM
o/qhcyKXDuVCfho1kCx5K3DTKATvBQ5z8auI3wis9KiPS2lTwwdPa/9L6fgfZzLsY5qwZ5dB4gOB
II2FRLrF5XK07oB5ixG7yLGlT7pnA6rU/cctzGIakGwHbsMIi1LS9etfLhE4fHB7ktBZRs3OgOqq
PSR+nLHBfux4F8nvfAjh61tXraA6APL+qaHb61I4o3n1vl6y4lEMuFP5DN5LUzj3+03yYBRRDiZB
6xvSTiboB76fJVSxluiJuzCzFq5LywOSmPnK4EHlCv0GxodkavhOJ5cJJ1GJWDi8Xu4sMXUW9uZ6
2xukspssZQ5GlPok3h1rGvbDIW1D6tfErV9mOVYrGuVD5ZdCrPy5aJjVZvE+o9Uv0vNqCvGPVRZX
Wa3rKk5BM5CICgOva948NpEwBRXxbX3confm+BK+N/qJZ/4P1wHcyV55icZgRfXsN59bEkA1QI+0
yUUNmzxinQR0YSFrEQXlvEU6eLcQsC95hUPpiUREmP/QV5m3SuXdVPNw00sqWm+CFdlOrClloRpo
qqsB2MgEh+uhUK9PG6rlb9gz+uwY4ZoOO6JtLNzjx5Q74kT0Mc3dzzT33LXpdCGAUwS78jwyQEbr
hVcW6OxHNcMUdnYiBGZr8v7gtc+aC594oasqHiSeYPvETp41WVICuGgOiKy5EvovXMC7EKcK1yZE
tFQh1Utx82RFJznztYR58x06MCUGOw8lhkWcfGu3Vk19k5ovd3i5MHymz3pMX/dkX47rqqux7UGC
VuzcjY1nBNfSb7/vCkRZnh4g1aIqTJwHXrAGM0TrzvVn3IbSsKBGBs7+nWRVyAEiAXggtooHke2f
1CQkOd9L+ineqFaIF0GpV5vb8zHzlYA35M5/MZhmgd6WSJ+NCM4aA5r9kgjBYyfKuxVu/icaXSJ7
kW8ZTSnhWEJ293qO8sYS3ATS3UDMuC91Vh/zxCvEkMnDVPWZzSV0PMZZCxCNrIpm67mHIrWewv70
GyblB5l6d3kdjtZD8M8CmMKVKUUiLWEQlAzGe90TcOpiBZX27Fu5wLRjXjvqBeuEsLy/M2XI8X+0
ZhA8Ckdr2qi3bQIhJYQ4NJhBvQ+bzDFqnh8dNEiVAUNJFcQit9GxLDcM/oCh5npWMImBSkNNPAFt
J+NTv8hMXcMNopktiOeUGqZp4//Lwt4m6LYooJl8FkPJ9Y7mKOrHQuK8IT3ZKMJb5+G0lKLaoC2d
/OCUKPo/5/4XxAfG+TQ+rnVjaqdmYKjezK2tPj/rRn7MkfyMlK1cGTY2Y3+M3N42izJ7mIBvKA6r
MqIKsXhhwO6y9wgoKh7E20xrOuBQc+g64+KzPU05dY49HaXmNdUdJRUaBVJbiiBdj06AmG8dTgDh
rIqSR8HfRsLVRVA314S6j8fMFFoeZSFGlDv4FTFCIXDzkZ+sv066a5n23QI/v7rodHLh6NGw5YAu
cObHPvvdAm8c+tRIgRXbFls4ejNGfwhqARZ9FUwi/IUwbiiIriULrQx97WJLAPUqg+VIkgvixgFC
b7ZK/y/ZnNAq/70Ff9CgKs438kVo3S/7FBSMLy8Q0JaCeV4nh8didxrc4SxrcZy5PIibZZziUl7w
cmW6Y2jiOwGIEow4uKxNQfSseN/I30aDJ9062gZLnWDI9ezb52xUHBEaZDgtjyw3qj3ffqtrlPF8
MnoG0B+vwunFOZgVZhGcmGMr8svWIV51mvJ2AJvllUW2leEMDodcAWIvhh4B01oJ7+yh4ORqoc3J
i4Ke/vMoQmm4otMrNngjrvJvvNLKeD87R2GkZ+uJdAsLJiFnyL+armqw2IUFnOjSy3Cw2aUyx5v8
H84NFfh7h+EfNacQtkfj0zQpGw7Nv7gS8rRbnkWJzoW4te1SobpQg22ptxtQXowa+3oSvF97Fhej
TokXHYaMayQjsWPSMnMmNmreVbkNzl17wXGbEwWShfk1jwO/DBBOgFBSmFsWInTGjJUFkPcjk3Wv
IOR4KIfTsgUmKF1OW0m2NxUNRSqX3GkYJheUeKEYhVbFk+515sesYsxJ0upnuZC4W0Uea+Rd9CkR
Dpd7F3WyZ7i0H+PTfkNDkAeSCgS4A5FeNe3TAFeeg6L5V+Z3iyrdYx27jUl8oTMpYbpH5deGO4Ks
PuxyX1pxRbP+PhA0+/UqgZPQqijJeZOYMtipyljwuVetBfLq90+4wlO62uSe3H44tRHNpmH+PkDB
F9hjVaGUTIHagLNaqItW9bMs006b53N0cmyfeN73fjrjYbUmjdldOJdylnfo1I6576DDuGT60jhY
FE6/FcCbgP8rrFSETQdYrGsb8qI1Lp3dtbupn8Dx8U1Cxf1vAFVUIfNMAySwHsdeKm5CTOXSUKBb
8QOAtIbwq6iNxCC0CicGF5I5XDFsoVeq4Wkvobp45pYCH6PCObQOwcAbrdqZMRvuYnpN8VXi8+Z2
VwZDXMTWjnnfTQsGHBFV2KrFJVZMgamDlncSzY+GBqliD2L5FIVnf3Kpknj2H2Ur4pic+46x27kq
rdfi3hT/SZPt8qnDF7vGxYOG9RjcjH28qSPqWSEKjumLRNozIK/ke+LHj15cngjZVOK3S2kSMXBL
7RUgpLtKX2ktr83EZjUikHjjgrxKZV/8X6LreQThJaYXevSDs+jHgrUyE91gwswbtIscX0kYyP0q
n/v9d5RKCTtH6dCkIuyIoPmR+91+OEYRfLLDd4d2H5mLmZZdkzbcCHHb/hh3c844MImvdFmkzA8+
i3CLx6TDczoaIFZll0DC6hgP/6/KuUjsF+TpLeQ2YncYwOznOAu01aXp/Fyt7mCLniV5GRVwM0v8
PkrOnHtiCwLAuUll64q75lbMG+jxhRgodY4C55aKHpDGTyL/4RDjXk5GQFNSqR1BX8jXiTUmnwB8
BvkzKqwSlhWrxydYCUVwz2i7Jc885KANcaa9T2H7qsE+trrW67YVCNL07kCssmsDQ4jgeFIIbpsN
ZcJW0tXJ1jThcHcot69nZ4ZoD+Fd3xOmKrsZ8DFg23z4BhrdKA1O1B3gsYlu35zlBkgXCD/W7yX2
jnaLY8iiMF+s5W6wj1Bnwh4LbvwWgP5guyW9FiDRGC6NZuweE0m3oOENqBqjGUqXFVgjwSpLX9We
RmT1Karuz5zATkpZ0KMZBwRXUgBZI8249buhNs8NV/xeuOSnos+x3fgMd1CGHrVuyjJjgtCqrqSk
J3xdya7wJ+GfQDvGcstZCHr7B/MIfqARGCq/IMIi60L3oqxNRm6QhlSbOR8la3yg/ZR1UoRSVfTm
NTJpaZ6QpOVk9vLMqcm/ZdxtneNKKe9VqwVU76oUBnD+iyUKf2wZsl71Mbo9aH2wWkQNHM7PdKOz
dC4pu04kXBZlNhuK/cOX4r/X72QNbzCVROfFEQCLw5EmER+UZtjnaliEdywX80Mtg++bxjXFk4ro
3LjJHM2sFC9wbp4jKgQeOn6+ou+ZoS5BY5XF65noHlOyvZVHEf8nOuIhf+Dm/gqHmKjm2+5v6WJk
mN5yB+yy7PQj2f5mdw05CDQG+SrLQDynyhEyyRT+pzdui67kdvB7BclHTmaO4SXJ7i09RN2fVuxW
qSN4GZt6dyDBDDeK/W8D6oc/ImyLfKdGBBp0D1J8pdwk5O0a20uCQkNB4QmpiC2p9kecqWYVXRzk
+ZCxTM2thtcsMi+MxZL6YkiZr3Q3jYUYhU4JF8xj8PrEkBIEqCTBPDukBaP/NNQluCrlk+uMmOQY
KFXy2GG+bKD1QAt2llFBhtGsW6fLyiRB8SbzF0grRy8dsWVbLXIreD601N6uhAIK0EfHAR21YoFG
tY2xALZt3deOGGNvSAPxS2dadmZqzKFSU/XssUB2M4vhTnOiPAcmN7wur3QffmkTgzJWBXRywjoB
SwmiMvYMFFiCdH8vmtSWD++xCjJeQ+AEoEkJpxYn3JQDVdc02JUqaP5TSPCDFWB+RnEzkCgitMBb
Fe18FX709/7i0cwroHTN9aH+4V7kMgp7yW4pF9OAqh/AzAMofIHUruMoS45w+Rlf4NS+z11aZYTT
QOxjLQILwTKFbppCaHsvDai8H2buVlJSzYqNFTxhedwoBPH/8LXS+dF10mLjkDlthmCQXuTKaLsy
CxXkqek5EO0zmsCQ/CRxjbhbkwFO5vkg0cRRjGzk2ED+WUzyEhInITFy9bBbQmnKC+FGtH2JRuFR
15S/GcmLjwiVPch1VSDjrC/UWD2TZnydhOo8KF0UHCP7xag1WIQUj5Ol3P+Lms2j4Ifb8gMzzfy4
74Y/uRZvSxHF2nW2d9VTH+MN0GQ02GrYDnJ2p4P49RCMcArkoD3iUWVtMHt4KfpdTLTVrA4ZMDFH
hBEPOrBw1VlXNSdz1fDwBdbRP6yRvVCM4IqqkWxwvb8LYX6cch1W99Un+28u3I2sMWN57Mcrorxf
YttSlf8UoNh+ugRJaK0Gp/y13ElHKuv7FDKIkP6t9+TqzAAfn+6++L3gtAuo8Bt9e1+pX0ArmMM2
LLXKA6yx1884byUu3uUEXpH1YYX1nq6sgZfTgK8aYbrOTpd3aEQotk1BSonhX2838/lzd2jimvhu
JIWLFqU/4qETYiHjTD2K7UwGpIUozUGaPCobJbkJfpO+4PEOu/5+uJfGmGqzOkaUGO6Fr9fhE9p0
d7YJKHOvi5UXfogj4QLkGBYo/qxpYrh5ehJ0Lywep8UwVyA+X5jYkpqRnayU3rumNhDMutYmz6Y0
dxbUNjfU6qGW2CS3Riap5HrGQCbj0hzZYuOCFWyWpzGzrF/KXLtlO7QIqn3f+nkW3AroUas+d+hG
0NYoEIGGn0ouwi22Q6t/x5XukYvWkUQA9QovOH27qcRRNJtDRnUXctMFhlrs3vNPKDEyhbUf+DCG
XPldh1GKLc4y4RK1MtyANE0S4GUFD+gqEQphTTgjroKvBcKrXsVjif73Xrn1EhmZGKnFfxYG9UQ9
cPWERYIRFXO7p+tzwa/a62nzEyv/k7SZ25jwgNxWr1BDlIDtdpfnBS9luNlTQtgxH5ZqgTJp+RWC
o1MsskQZGXs0XjRv/eyHSGZKCKmj+ZKEz52zkC2khdOqW9PfS/RZ3UcH7zcp5yPL67S74+hiJf9J
KOy0e6G1NQFCFgUdNjLHo7Z3xTpZMFvkhZHWC3tTVLOOiRbkfWAdcr1/2GRtUbTWSirYGTp+YRU+
9Ergxhhm6UBqVnBVFtNlAKpXhDmtGtgsgkNDGM58cpBtabR34BbBF5QyN/VIRe0PMYm9tj3nNaFA
ftBti5rTUmOzutma8AhcyjWez/9Fj7XhRDNNWzXzsLwJdPjc7cYTYTwJU8D+GbnYeQaLZZTh5LSO
G7O/022/OYhTNjPswM15Au1GY7seT/uOHPr6HqCfoQTyHul4HKFTP0SfpYIEJBtwXEoiGktxxr7S
stj52TnvGjWw/XkUpa5u5+p8ttC109lN0zG8FQlpyAyxt30RjFf0o8iNP3A/BjllTHX5VoAiajRG
XLfvbCjkxUW5ZJc95S1dt2mobVa1nin2hXx1QGpvhw9URf5UWTjYbgTQi+Ze+vopi/jDVpzoFOCY
kClA9JBTOuCEH/ACIwcKDI2HvfME+0INpldPWSs0hDtCVuEc83HQnnK2UhDn+LrPVXhqJhUd+Boo
g4zzj/zb3n3HoXJJXki04IDAmq/GTlFzb5gRrOJZMhODzKOnsEB1n8Oxq60GqDlec12KE5P0PIGo
iOsP8+bzcl+p2Xy6EhYA8x1P28d5BzclrTLicaGd59tQBsQV97lCH/evhdBFdaJpEzqFhKr5yFX6
y6lHUlCp7PjF8OKTLCxrmYCEjSfj/JlfOgf8FLcHBjwM/sXhpsdKEgxeEoNwL4LcAenQDfc+n/J+
vkdbREKY5X22eHbyle8tHAbT2J9EAPoRm+inuZW2bwojz2ezlD71Zov45/a+CtwKcp/mEySPZ26b
Xz5jtMo29/bLQVnb7Q3hOq/uTs5EOG9iQuQAmyaTDZrGbtUxxatIcAXeX/8eWdRcpx5xG/3I1CAX
0535g0oLEZFiv89CZEVywWaNunPoiSSJe7JIuj1KODqV7+oK/h0A5qUJeOXG7MRcTez3Ly62BpiK
XaAYruF9QxgH/IOW61vzMK+L/CKo9qD6E1dB5hJB90AgS1zpQelk6kGPyS3UR3XAWba/I8ayo/0v
d5qVTtDDSeTADGmQJk29FKM20Dgz+Spr5x6NYeKSxrRMo7uzuwqOOjbWWAeTxxMACsvtru4R4Nhx
TWFOSfBfjo/5HyhD23HKdsUlWH3G6DZV6CfhUwAK2xrY66EmPJJP7/okkBWA9rggSW/hGpALxm1c
C2PAey37jIV6M864e8SSGMnK0oso5Jc9GvF67Jy699oGok3ItzFXrOYoFigFx0pKwN2UIfNNToGp
/lb4Eyr+3I1U76jozSKf0WX3himX5HWaNr4H6xBg6AG9mSr2h4D15FsTeD27FAJiKeB/U/27A1wi
Cd7P14G2pyH2fn9Gq8uohDH/NtIfHzKT6HzpwrzVc7AZHkBoRAHOWO2GgoXbEPskgUpG1y1qbkyj
ASJhHwLf3dAFb75RAv8ihuT8YfuLHchhDmtJ7Hi2NoJGFelIZ0gq3qsiQwXWL0FAwkr26jw7g/Pm
6B/zWlqMc3PoJk2lByT+7umV+tYTJpjmkCmI9I6h7/J6Y6iCHB2C+boUsnAfftoJLzPopG7L5K0q
n9mllbCaID3nRzIICrtdDJt6ZvxqmJp6yN0M7FEfCMQaJGZ35a/mDkIqKischb995jUbLyix2vw9
6+KvjZkozSPaa+yp5TzrKAV2orDBw72LTz4L0u1rMO9gRZukWNN8hZOc1CbRA1VRuPE+CTU8zsL7
2JaoNr1rrpNf1IEaLI+P3a91tMm1UL0Bwd228HgFoWZbCMFhdnPO1jJL81moxWYfTtgTzMRgqPkY
d9ageA1HEAtMHHr0GVxM1ndGy0yZdWdvCm0UHmVIK4pc+a/JsW9nOpbbonUphLfMrtD2jepMyLTd
Xpu+TBMbCGXHaFkwRZyovKklzYykyLwX2g12zRdrsh7dprpA0F4rTfwcUxMoozs4fje/s8ZkItir
qYAEpVj7bPT+jTIQEUfq7n2xqKhISzEhUWvbiOUiaGLsv6jSFTLAqkmJzd1AFgvW/AWv6dpnxgZO
KmoCsiwuRrQ9h8yEFmsOTiG06G+DhsWgQvH6lfareAi91ihOmOYSgJyzSsU6mz3m/n2cHjyFNaTM
nkJoo/mDnLH7nrMwhyxfWX2CUYETEmqYw9XVIreHuMNPhWs5/zG/qEE873LRhJFpa6As6z6n9Jp4
BqhijJD19dK4LoONwtQ8lwaOuSIacWpg8uav/fCTAEbz54HHgmy3B+ySqkjKfQ3jSQQzrbfUs7o0
pJ5Ga4pHjoRuYrQ+wIBqUhDVG2ArLYUXDA6iCGTWX/+ihXKUaK92k9Yde/vuWVD7p/07cjzRziNn
jfF4aZivB4nv7gEN0Jhxfk/sJ+6/y33GYr/WGurVLARLx/XteTvaihqvf95zAjORjumFqWf5szM+
ENaCsh/OpbK/KsQRB2mSr7VWVwgTbKpDKR+hs8atUuxz1q2lKINTjl4uFZmJEpACRulQr6nS1Gv7
1DGHJPolGuQurEBIVs3Lm2rmcXWU2F3q/JMHuYFi42iPSy+H1MOgXlJdGppqktWAWTkv63le6vVU
2VmwbO9roBkexnDxC28gWTn5PlinbUIgvhDU1WnE61ZkVv85VmYCYbi5GrPscg5Qw2qfpz99DeWP
qmow5sHT0hBoEN5L46bPVvKtjRXx7Qd5BIqCXUYKheW50C4h561XNmFNSp3KF4zUePRa6ZrwPoav
f17JKcRnM2+Ey5TvzApzM4Nn+WsLyf/BYMhtYWnAJlZ2ogEI+TJEAGhjyYg71lnPOh/MX73yGg7Y
tECMT/5+fFMshFhVt+70wXyE+EN8MJvAulqO+p3QLnjmSLwJBEnu7aWtPAubxXxvsArxMOPcR+e3
4dnAPws/TjTGhMlLAsaD27kWNG5omXyLYOPEe3pU2/Rp+CVeDTDhUNPKaqrrLGR9bKIUQIVwNWhs
edrIAb4wzN4Yeg3plF1xuwU7O4y6SEeipXGE/oESIKkpTfy8t1q19HbPDROw3OkTpMjKBxczUuAW
IX3CKOQD6WB8Nnx6dydquHMoHFINB9IDxTGg/3UQAzA7sq1ISgPRM8kLkwP9suWuqMEA6z6oFJcs
a2mhb1MPDlsTnSjzw3WsKKpnwaxsVdCLFyW65dhBHo4have0s/YQ35E6YiB9wG1VZgzC39oqDB7y
efZxSi+s9QLZ/mSbVd34ZvKy91rL8eySLfNH8B2whLg26F7wggtqoBYd8BAatBK1RMW2lvliiD0L
N+AnjAn9evHVzzVK8WnOW0MB15xD74oyBkUCuFzyNYMK8S0jblATRvHXF7o70FrVXUP0qjskvzZV
236vY0mHdTj7aNuQqPylusCLpDANl+e2jHgiN7potMIYRJm6gg58yEDZhaxZguyybmOYpwU4b2RA
21AjEc1pk1VetprtSP9Qbie7oB7K+KvKqu8ZMRIRb/bRBegvltjYIYZApdm0OfPLqHBoKlqfJm5P
VirtOY7fBZxr3MuPcKyAjF9VGObCv14Rob6GP6FuWcaBob1R1AaISnNaEK0uBDxUso1K4mV721X3
1uCGz5pzI4zrG8Gqr1SFi9nKe+dmLr0BVXSAm/W8iGonYnWdQt+6h/Q8fgzDNW0ffuwM1orrf8XJ
NJL3mOGN290GVYpI+kGOB/mFOQ9U7EhYjE9MzBs7AG6TxbkUndqM8jz6bVF0vuserVxPzxmbU6Vo
IMAgEoZjIx2U7iQz4v04Yk+XX4jrivg96ZcOSEq9dzQiUJg6/FEhoxC8SZQmJ72EgMWYaB8+QvTn
XVRBQ4XTzKUEVIeea0HAm7A95EqjTsH8lXhg1dvIsK/P91WKNkueLyWJAnkscS3nwUR09n6LH8T5
T+SARa11TquHZFLTWjXtsKGtRqgGyznsErVk1PhRVs/Z5LPxbfPbvyzJ1dOM/U49qtxM1Xd5IGFV
uxBmbxCT01kbKCjApmgo8tZgdIXAGqjKpBiXdzXcq2plo5NEa1MKJNqH5z7j+p3lVCWA7bexkHQd
pPHny11frhVVBZasCG7JTg3kI1DG5eIIARqIFD5Y6sk4ejC0f19q9t7wGCjgWemhwGPJUx6XnO6U
UO6nFAaKlsZftBa2HW1X/BjnCBvssn3DjRMkv9xRIvvKVtNXmX9x4DZ4DbkxBLtb1UxC//cV2mZD
APPc/ee25frP1/saz6LnnnjhVb8PKk5TIw4ds7GAw0PLz06j6eflNmLSkJktbr1jIMjNSHpLdzRW
n+BkO78cb3AbCwOJT5LhxgKDXNK7VHEMoAJArxmM2y+L61pgpaGf9FmoGikXuVxU+lKef5jUyvOi
lkwWnuXGeruABnd/+yyv9p7zhsCRtmtQO87t1OrioZ89uIgN5rp376cMI61Cj5/RvSygI4ELPO8p
5ruzGy62fYPeu/F0wQFepbsTA0+SZWYJQHx2zN26na9ZlTFFjQ2Hrv90AEPc2BAHAAO3MPV7lGzR
u/U5mi9k9nFtHcztTX/oJxb9Im17NicM3yeRuzMO2dmKFCGrXfdrDxH7CGZIp0Ij8S859WBC//Xp
e+FuzJTwwJD1p0uqi2eb2wUdcvYct5v568z7VwFpV6ePufsBtuHYaAov3p6yPeAIbvt9GWYYqqPC
g0BAflHvoAsjE4YQ89h3iH+yZjL1Mj3UsL0iXEuHH9QXMSskVsbD34rCNRSszAnawBSko2zBnBYH
Y03V9bnfuX3hUrcGyyUcQRYbwD7Kvfm35gJcH4QpWMdRUwRRkHXyyeSYsqATFq4LB2A64ahqlXcz
PP7D0QSYHpoJ/yjC6CqlZNPJI545X+Y6sPXqPs4/rwiXvtBUh7XZkSKm+iakSB+3Yl1eLyuyEh3r
D7T789QdqqWd1T+cPqw2wZBrdmoQqRRncv9HAIbX5XEeLQYGRpPE7nihT9hCNFMozlgqABJe751V
Crl5Txq93/0u/a82SKHNY3cicDNbNfhmEJc2EOuYVxr+/U3+k0/M67oc3cCjusI8xkZ4CCNiVgCJ
o/3qL929r0SfliGeF1lV10/SEvtIrL5dkwyesuqWD0WnlpAT514K2A1Q/OTDZfyL4CoCp/HIQgl0
B+hH/kItz5t8sNeYN4i8dyuVXVKb0RyOegmmaRXwZ7VoCMAxQjQ1I9zqG8VW55IkFvUWL9Q2fgvn
jG2RaKuCi3bROvdVxsp6Mt9NOqY2Ot9fu6tn+JEL4ylQ4ko0ugNnfw+HyR2BRrS8eezS+ngEEgWr
SfPyYer0s7HMb1/gP5l8zQKajujKmp5Jpkymtxf/r5BQMV3AnB7BghQabdFaQuTP5GibEKnqnu13
B86UGK1pJYZKitQrk2/XgzHdExX4ZI08E7+9VxDG3gXOai5hqGQeuNsnzJ5PVOS4zPA6EmNbpQRy
RbruG2t1kjc+ZnFHQbrKBB8MF9U2rESZpcUG0vix49ze6/sNi6nZ8xYqRV2RhRHQelnnW8BXjnL8
wImpajbN2Gg6KkadvzjMYR7LNpUKO9pwxpbKAZ1g1QwzUl6jG+nzW1t6R+PZBvyjqOGZRena2GNx
V/8LgaLU8c0ZDOlr6To+vTUZnDvnhcbe1Tl5dHBCEGapU2FID1yMlKPGYAOOi2bkSPjTkXhyapUA
SSZeFLZuaYBjJdwu6iavcTs2KLaeYKDwrMUjnvqPPyDQZQd8wjcfdOL8LEvyOt97asAFxWyVHuKP
SL9oq5S8P7nLD5kwnrHgjfDWUlHhnEYvKYRgTUrZ+zSlVroC26Q4SWipzn1LVrA6qpNFLF+E37Y8
g3KmJmVoSWRWW2WOeW/ucu9K9XBgJpc1MeRR0sAT5Vc8cOZsL+lU2InPwrLiD+7q24B+79fSUxFG
uyLYDs5zweDrVU3KANkk7J6n76HKa+G3izgr2iUFEqH00rYoxIvtLY3F4hWcnWUeIfl86QUHyX1b
dDP6KvHkuEg4XuK+QcZnSM+KMJNcxu8AiIJJ5QST3p6vkPrYUEgeP+1tkwaaGvrnoy0A/EgKKR4Z
KWcNvGH4WptI9R3NE2l+hqLBA2I2yWpDIHF8BPhoslGdbOptw6OgukDRAI/betN26h3A/zIlmOZc
/7FoJdNOYeD5vXQC7RM7k/GSfi8Iv5l8i+LKdtZBr8oo5n54hVmHor00tw+KiFN8B+RmootvlYxk
jtrh75r9BjFXsWhROkTi4Lp4oUY2y2FsKOlCkTgS1CyAdpjhequxeV+u6qjC07V6wUicVI50kCjU
mHg8OJORRKL67OIYd5PawRchYMSllwdNQOFV7vLvRz/9GBL5q5eY/Wmc9XrEUR+sCM101M+TVqnB
hyvoIPrLTAjskLfwGn37L3aTJUpOvkhTvczq3bAcKjx60VY2aqxoT3QZIOMxOJwdPCX6zjrinfOf
obC9xdzcQPDJmed8c/kpY+0hS7HnZ6VcsG8WnFxSrl5ttJ64st9SJ7x1CEqTZjUIAC0GtM9+U47i
SnUBgg5TL56mzAiRHFBBNVO0FUqc5uTaCBOmT5Jvind5BUXav08ME+iBLe3he+LSVrP64RZFEKDf
pEFlS/l/DXy1Am6sMIkR3SAqgr7ImVEpbgN45SLCex4CN7Eg9bbgnuHHbQQqHUA3vvdj4aakX4hZ
QCMAQpe9SRC4u6zahlx+R9eLuS9xr/BKxUjUEahtWKOeO5UAjA78wDr/6Pkb/LDFYoSip9ECjHB+
904YOyFY13+D5DN1Kt37gG5YCKr694WOZlva9FS2U+TyS72kd0ExIP3KjaqbyWiK5LpPLJBytUrj
QtM4q5aZr9fGCzr3KnEZEdUYZE/ZppAPkqbkTM2e3HZLA2yGQzdkEe28gaQncZVqyXDONWg8Tatn
oValBRBLyn55lopkmNzDG6uiCzQMSWzAkSY8hNksLIS3hmX5OOSyv42R7a9zGEB/t5V/9PC6+Z4h
67zdP6hoahDOIRO6nltV8wviYUIaptnImmvfSTxPeL7tIz9IGxBHmxTpMFqA6+jgp0PM2sLxFlIZ
3D1XlRndPuV3LWaL7YuSGhSgmVZFcTA6PO2ySWCbCUgfnt7kYRxYUL9b/VOHqmZOoRUeDDZ0/SHi
oEDFKfwMiPyuKpi7VgUsBAhJF79ToLgx/Y82LDBZCJypMcdHRElmv1TkgDpnYuZ+0Vqrj/dwQ7bE
utJl2Nj+3E56OUYpNzmVttL1jgvM4pVFIPZ4w1JUBwsjsSSTVa6P3qlf3kMi81bQVcwOp+a1Uw8r
AZv4/5yn3B7+0bqhZiRwTMbdrp+Nt/NDJidGh7g3zpVHxI0jBQPdGwVz7Wgkw1bo2hbEJjdHvKd0
sKGwqApyhzYg0pzVSZOs817VI4YzVXv0StP8CvFmAKkK4Y0UaSbauriQwF5D+GddXEKJQhkjSCLD
s0xWTlX+RnOqGbUQIU5VpR95DMtFwidphHpiEPur4oVgZwY1dgpk0hrx1fkVKr1iCuqs9hEJrjKD
cFV4wh9crqLB47XOMBlYAy7wen/Lglo7fs4i+EYU1k1BNg1ZyznTjHdta+RDk+kgzcti2VHKyZSw
sinlTR+s60HUwHPTrkClHOMHDbKGJUwOn/pI+zP7bMIy/NCadtLLu7+SvKSxUNf2CmpHtmg+IBsm
nuZgCuM5mxuT2v7oJkPIXf2McDPBAQqInCMttRTH9ffID9PuZKJB+TGnjaHMOXKel/Ixgicjqwdh
WHbcNI7TTPTesJgvaRV7cmaQV84Zxkeh3gMlDAMMv/nSyroipqkPOym2fBuEKTpt2OiAutA1iD4p
rK8TWA79uAwY0+dKvkYefTsATBWN32jC0msZGBZD7MoLuugeAsNKNg722lNlnHHCodGBcn7fNlkU
Fg3aoGSfBqsB7JamcaAn4bPN/ai61TGFO7ZsQJ6Uhfpx7tv3zvvaYLS8t+Fz77hoQOVyKhu12iyE
pY3DiPeow/wWKDzddcar95B8W3x/rmadhvjO4mKFzRbrp2/22I62E1XpVTOKakMuCINjU/Gq2uao
Q+j3aowGfiaIMIMbDAylnr5j4AJOjhJ8zaoNi1Jty8MKusg0cx2VLBr8ntNSZDILG5SOog3GxHnQ
iF27GkUSSvIwZ1IbYZrRRdAafZynaPXJ2HLfYaxJAb3NBJ9Cx9AUBQn5mJL0fcqYlyhdNizRaoN4
V1kQ2y5EEOgtLaKqv0dEvbokHZdN2+ak19QHGaWbEMd4A5PwSGq1AFtYhok4dI2sdYatdoAzFtYs
G65wczXc+1wKJ2j1z5nYyIqNreqnVK8Fb0GSa4RK/wc3yOlq9DyJQrvHh712oVOnVfITyBADgX0Y
MOpmeGcJSa1Zc41Dcx74Sog0zLpMedb3JJDqJwIQYyTNBeDOvY+XQbGcSjX24ULSSDzYNO+AgY5l
CjdqsU5IlvtRbIh1pd+4Tt/+fHGSaH5D0N4MV+ALMc/uc9udOrG+zH0GnM8qzMSuAwkHouXFDbL4
RPMFJzqMfWRH34yScA+japzUQ3IAEVzCvzNDl/+o/vLYDteUakl/PaMKlkqiWDDElcdqodLeAo0B
sj8m/UpfXNw/GQkAQfHplFQATC1FxZZ1cu0Rnp9wKjgzbGMuD5koyqgyhT/cZbxuHINIZ+aLD8Or
ym5wfOQqZUicExNNibc8QstWzwxu7ChY80DoeJfc4VKG15rd944NFwgWWTgJblWqUA+unMnqkZC7
5ntu26XGH3LRoSC2ovMXFaHJA0/ZIcVLnHVh+v63QyZ1Pb7gnTQg1ejUKLLIC99CqHQWjZ9RqUlO
TJuCs7+s50mYc23YSZMYeucZaU5l4ldwxJuGRz+Qjes9TZvxtI8qd+ER7X8qx6aagmCmPHXO5/g3
HUZTDrZKxifUaKJeSToVNk3lk8X1hGOI7Wn7Z0iOOiw2F5Lm0g9UQdsaVd3efTEvI5wWidCgk30n
CL5s7elYVdLSon1n2xqFsfVOR4NpNKFq803xw/Z2JWONfIbpuLdEsZvwAX8PnMBO39VfvtjzeYul
tfZyAvVyM6VlF80yQOBVY4jKvzfy+i30dB0hXHAOrTbKX+Ku+MZbcHwITGqwjKvzV57BhhlL6jK4
U10O21H5KbPHvGAlIxNuCBxvSO0wsiEAMGIsPulTjrExj+vMawL6Gt4yjas8vEWq8yhjdXKB4SLd
EqQoknewUG/MC5LSHDrBZPOCkx7VQktEJppGKUUfVL2aQCtRO5jIiSz6hnAimDKv8SWMuW/qPlLb
UTMtu3RdQsi10HFG7sw9Z6pdtVBJbMz4y9MVOs1PrCPN32g4sktN813Ew/xuM//4oc+8eNLei1yt
d2lVGMDR1eYjqCJInxxBhwuzd/YOMpJGTKjdD+KTE7Cl82T8T3DLRM/G+iEfsW4ieRJYQ570IzQ/
qKEbgbNwQhRGDkNulCv1LgJCXsiWM+yG0tQNGEh9FSR84RLHoiwCRm89UdnxdYwLSejZAarbg+7W
Q1wXa5NCr0yWobwk5i4d4+Luh6cdAtVCWlnlUgaRK3fvCn9EZUChm4agY9qJ29JCwwdrnC5ThKXB
DvV+KZJT/7RWt2/YMIdivvagrepW02TZFYImQ1fEHUnlvSo1UiRQzsx/cwqRTXPSx4Ae4Mq2YICg
DI84WjEDYV5BeaglIHLj76OlAkeM9H5NWhQLoA04eZ8JxFbmvCjvksjoM/fZVk6y18R+Ln7LVLfz
XmnnDJjYVTjq2gFiGHzuV2JbQtEkNPNWux1Ukq53cv0JO8Dl7PhIg0sLVhIUB4vgpW7IVodE0aDG
wz7GGeYhhUwZTi64We49kuVkpPavEQOKZwOfyE1s2HJB6AeMfT0AIo5/yMNW9atv3diyUBc0TAj5
cmi6utAFtoO/8G25tVxyrzZ5CEa5zXErXhm1rHKvX0WTPB5+I0iEmMpsG+7ubqitCAVKhOKMEviY
bdyNOMonGS6K5kuJ0HhjuZMwvb1PR+o/GQqon0F5jDUJdlfpL9+cafhGf1BrnFK0w3DOYXDY5+zU
wHvxBs9c4LD10fSs4GJSBr6BgQ6dgWkDIURaSthHV7Ct7ZW7/tcJjFEXI32qKTSrfH9v+JK/PEHV
r2U1WGhXnAwYQJP7J1S/cwvMOIvIaVYL5hFarSUO0VhA5MgJ8S/azmmKENVa9oMS1/qTYp1wulG9
6DA1zsdK4wr+C0ckgaQbL1BGVKilZk914tmjOA1RQxmuEadtn0dA83nePLVAP4Xaey2ixl1HNtAI
HpWcIbMcAodyoGkx+Z0Iyou5IroZDQMcc1YuN5Gq0c8xIog+m7iFx47kUSy1OSszkdzdt0Ji2RXT
TENm2I3jbrxaoEWgQTjm4GKAc0ODyM1SsCAjNqbYSbXwS6m2ubCuyPBaXxVxSJ6nhdsTrI8t0/6X
xHZXAOP1fGUXsA2SMmvJPZcOsCyu3ipqGqDWGO+BWmpra+lSykyS3T1ZnL0t2Fll7Bq0mLmm/B+d
pOpwPbBZqL2r2D0Hw71q/smHfYKrehthZxJwx7VbHPo933Sg+g5Bdii+AuvmauFP82rPAbxNBQVF
HC+Hj5zNo15HBkycQs5AV5MXaPJuo1rcgzLR1pYEqj8K7VllGUlKkB9BZkC6/5lrKdf09YNX+Ou6
zktmTbgzsLXt93pbNlzg8bn0kR/w29TqqVXIzOniP/dy/CF0xTRZ2CM88X+rf25cIgYsdZCGnkAT
tqpLNZKvW75jdC9ekdfhGB43A0q/muYJw23et8EkXhGbsw1VPeF3UVYKh9a8+4GeCzEGndwYOwP9
R8PooAa2/p6cEwsZXvk+amux+1tz5hZ2dg5//P/1sO3XKjuMXtw0HSVeGX8OrzITM2xb8emseoPA
QNByc0c3YGC19KVUuLy9O2bWSkXzJk55nTR9SwQEVXDJaKHtoyaZwCRF7H/DOhyY8sW4uHKY3ZWi
IY7pG6fUPmhyU6PmaXW/Rb90Jt6joD1dE8Oy6ofpc7bpcIf3ghu2a4U9ZgYzlt6KpJ+LvI9M3AXS
c5AGPsR4i7CvUFw6+x4gffsas6d5/n40FOtLrgZ0R0PBwLCrASXNGWjQ2F8WsX+3a7/p4c/nbPSV
zopvXP4DmIrUyCXxeqPAHdZ1vBCTdEkxDM0bysze8vsEfflKFTtRVto+GjuY2RgpixMvxodG4pIW
se/eRfWbFIMsWRhcS4OMDp+uVpKuGzI7LplUM1NN4jyDGwwgfMBRsl02UhJXh+OKpBx+AWsgLPmw
UMsPidfmRjpGDHKi4x/+Wn9IoheQ1Y6RL0fMScT1H6vl07WraC4DBKfO5orADr8V5rMXqaV+lks9
y3WFh/fHvhq0e/+NIuSF6pXS2uAq1E9d9QWjZGMSIUKM9aI+9W4e3I8Y2scsINlXyQVZBtcInjg0
dAYijZ14f+9DbrijqTP1lCDmau2RO3DHdrAxHe+CDLc4p8SctnHCTKH+8Gl9chvjDUCgDnDdrChH
3nLi1rEDL0Gjq/+efbodpNLpy9+yRKKYZEiKxPvU5jOcdidy0HuDyy4Gm6AN54mgBhDTtM2eak1L
q3uptQYLvquq3OHJgTsbzQZ9JBjcYNx8PHl/EzmPqaT5WTRhwiGtW7Ndecl3a4Xi67tUgSUtqdGA
FXsenYG6L/AjwleFZRzWN2c70Dv56FfaCFSXfcvqaajsWtlce8T9QcIips/a6iiw5YeleOAwTLSJ
p4oAwjiIIMMSlrLbOxeoZfUyKfxFh27GBmHEN8vsmmPmEBEq0ydhGZJYvVFMYja6mexiDn5uSyoX
OBhvUH3JUlxK76k5piC35nR5JHAN9j7gFNpJAt2/hbeeWnFFc1CmbmYMDBUnKR+QIW901L/dpFZq
vDJ0H4TqypKuPrOXGHZUIVDWJAoR3aFndH4TCW6bOd6eNwNFbywYW/vb0LQDDxnk4t4jH7MkxkvJ
5T/WHlrDhgiV1LBc4qKK31ThPowNFSkp+mxqve7uk+toQ/C0KmXn7xYcCxgeoYH9yEH+kA2TP5HI
I7j6xtJpxp703OA36xTwvqnYUN1Uuswa68kqyZqx7G2aRynT4o/KCIvJgSzRQvVJjLAzSYhkHWNF
fEBFGF9ha6F4hMb+9Fr9am4Q3BHqRiTNo+u5A80+i8C1pME1cYQwbdAqaQ6AdhOPx7tj197CaeSr
EKsc9OBsN6sD6/f/YWdEiZMXq2/1Rc0+RRlWKjkS9XDABa6RCv+TRDlnotPpym+WgSBKLtnHxBmB
5YWr/no4HbLY/Nx3tHRsJzgHyd7oJhZf8z7taGoNOkrihey0053RjRwlnkHL+FqhyTXkofJ4SoCN
+aHhLzule5I5XHgPKJ710l+BvkV9B2Wt9T5JdcvQUawGj5UEMBpo+5S9+hol2lzaPbD4DlNLweJH
U+TlzhWMGI0+gP+zKeKzhwXTH/jQDehYDeQ8tNhfXVajYAD5AR6enLTQy8YCKbNreE+hOJ9+v4KW
ANEWDgwwkLWwXFX339Y68j4RE+SVZbQiMBKEKMJK82MWIA0wnZsEqzepbfxmWvw1qbJse3gfiR46
ywW7KHlmKAfy+0VmP+N6EJzKQgJwQkrnGfJ+xY65EHB2ZicL3yZs2UvsMslTTvVxktbUQPXPkEkP
yeHJxzA8CGvR/sygAfsdpr6BxcdH5hS5xhFiReesr7UyN4R78SBE9E96FyxP7x+2c28qmrg2AIkK
jcFONyu8jP5oYxDqCI66pWBn/0Kh3WluICgQA43P8Cm8bBVZWzH4w+8NXQEQpYSQAxQZrRbW5UaP
pjgER/6tbONROancxTI9/twYqAO2J39Eh9YsKtyMCBfwLkV2FZnPdw0fPmTxpbk37MhL2zCz4PdG
uvY4N3IHs14nraq239pc5jLGzu8jdqKfgcZPQHm/ns3Eet/9Ju8jcz2SzTwWk0d4DtvXHozTjmdM
T6oAv99HRSp9ygTwwayu3m5Od+8PiSkOh0QQA2Tmh1vc6aUfs388HPjGOYW9GYhtD9VEkDNxwZ4g
OGZxZJV0CBPX+qQ5n2KXW/qGyq3UbgyRcC4BFKYeClTOJp0twDOoVPAzkT4CwtZP8ls9l4romqry
+eQOHLy7FVCFjw0VvJWHyVxuMRHf7G37br2AHIeMk3Sq1kuiHaoi0ClNZC0rZn0OyK28GqzpT8yh
gHcliOD+BYGVSH/Kc1BPU9vqZMBvqybgn+TaDnsCLa6JkrT3vpi08ZdpL6XP+cU9BOlWRb8oV37P
YKeavgCfN/uoSBie4RRQcmUzfXxW3aaKmnNWoQ5y23Ak/KFCZBFS3TEJR39wrPBeXfq/XOrHCOr1
bRPDnrPO6XiLzNL8wAqMfpcPYaBnCa3JPFJO5EByXmGaVjCzM3vGa5LM6JW3Mx60xE4wqli6B/dU
F8XzSyYb5I0V2IU6UMLN7BwbaId4J2Z9CzLxNiOfYoX/6kg1N9Xbt5BL7OVpjXSbWXS/tqMoWodl
kc2h8NZ/V7CXjB2aX4jjaVnDKFPXOJYBxWCeHOBuCnxISvR4znGtJagDXemBswjp+lw5ezsR2ynK
o8eqAlHijRgBsrsNVLQESsDRiHvu/4tsYTzrH5AmBkY90RGpja9mMGqWORDP+PkcXv/Bj7ePS+Bh
IjvAAlO/o24/3QcHrTmaLnL/ztflJB4ScO7BEGfYh+p7kZCj4h3P62IaZkSPTOUc4MsGuR1ZhOmW
w15miITvN79sRJnZ6aYxWwMYfAGbw1wnKplfbSymZgEe0oSRCNm5qeKdzh3vwA8UBoVe/MXv0G/T
tNEfW+22yQTbTgeoofanirs8W9LF7iA454KDzQtLpBMLjO9ZuujfC4ml+7iqX+nITshN2pdr5CJI
9sLgiX9rt3LRAyJDmHJEtbcHcYC5l99IDl8i6yDKctcRPhpPSqEsaBmErRHvacSUH1JOzKZwqdgi
/obSRjJQzRZd5cIkq4K96aN5vFwGtDTLRaEQEkkK3BX9FAYI9c0cgjmiNCsp4dp100VNP2uYi+E5
+W7dgQuwYoRJP+V2YHzg1dzFRwSfYfMi45LV3tYAY7WlDy7kTuCb9M/G9j9y6a9uPy0dwjHopJdN
kkLMVA9S2HrQoW1g4muutYMdMjt1n8CDPI4K8vsuQ0Xd++WFbDt4oU1DVEp9wIFa6f6Zyq6uJro4
qnmRuFSq+931H9DoFRDthVBEgaC0UZnKE17bHSPFd7ZatOpAhoyTid5SHA150lFhyGEHa64hnW+w
D7Ns61BclSDYrduP7rg=
`pragma protect end_protected

