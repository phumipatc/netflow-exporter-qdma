`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
sJyx2gfifgnYXxmFxYSjQc/OS4nAFs2hYdS3eFe1vgd+evjmnLlQNfCzrRL00KyICRwryS3x0lSr
qHz6xWWSa0iPpong/RQ8jeWoZciS4fV1GASwvrldxBLfqnAZFAiZ9cMMqjMP0mEtFP6PLsGG57Qc
07FV8iAo2/2JQ/9OgVHsbSzgGiD6qdvsWy6T8Dm064oOfMABd60eCGRy3sPvoaTUYw0noPkDnzy/
DeFVKnSnf7dfPt2estZmaz3Duh2d+A0QwpN0Bsz9dRS/uN/nLE888fTAWg33+cno/TXqsRE8jvLL
3shuYaAIVid6qEsVAlr+9L4s3XlwN+Xrc9BjdQ==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
C3Y51hdd+MxlyYowQDqekzhMJ5KwR0IoNrpy3nkOqJDwAw75ZGRv87AtuaC5lApKTkBEg4h/aqsv
C3kTTjXPUjWm8Zp+R405fTSmYoHSnCoEK4AdPJgmLJXj/yQlZawGYcxCAuErnprPDdhaDNfGwm54
e8syXSH0L4Y6zq0Z41gFYnr0cKU10yb4KmHij0Z3WfFBG0o6hWOlfzkepJebTxgOO3uvWxJ8/Oqq
4MLV9EnIzRsp8bokS2JIo2y3AK6kaKAq3ab/sN4Yaf2LzH67uFNPafX5041syhSZoFIx7mL3wDOZ
UaZ/q2tny/AfGTUN4+TV5UUew6iQM3HWm6HL1wAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
IcH8WMm054kikAgAE5UXhsyLV9hQTGU4kMEgksLdrGbaKyLULWWmwwOTAuosIB43E6NONmfr+LzZ
rbKp4l+CBA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
PlYirIIM/iseuaLv4aISkQQhm+XLiITTLDM+EGloNN+0y3tf0V7eudjnAu3DP7XF9s4WtHv60rZh
ZMNmxd8X93UBU+BFB/uKN61H3m1TQMcn/mmBFYiibciGMWuv4D4UAvdRciWyguJyjM05g8ucfFcb
Ql0cmbM8j390AWroSoPo5vW9ETYYSS2MPa9kP/08ZCudMd9+SKPRYVHKPHBVH6ngEkCrYYwsnVK8
AIxtInFSeXyIH7SpwZpLglElcj1pb2j97Yh/T48SC1ujmzN88H5+sFnxoy5OiGSrlqzowPzGqPn6
CDQWS6WdwNH1O+15LVGHcjgV5YxsuIMMMOi+sA==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
iXzGK+MtoOLqjssfsGugVtRYN8PGz4xeyVsrz4u+W8rtuARauCjOpgkWM7YKBp5ferP9w1o55Azf
wA4S29lUkW5ESW9Jpl2U4/oEssAeZrz5d66QrQDr6qG+Cm7UytArUNE4O9/CeDlTpr2seek97LPQ
iaOnVVOk2UWcNLUxnxwPRcc0vk3YCI2RrbAnOGx4aV1097SctNzyx3EQU8Gj7twL9f1xIop63BOk
Wpnfi7FXI4w5b30HTgNecMr8ZIYfxPYGMtuGRR+UZb1AjZ0D/eWH1kdPDr1Ln+6V54Er1ZOUnwce
Nxe677tF5C8yMWcRLz9JMfSTv1DtOjz9XWvAUQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ao/kFPSIqDU057oeaAzk40xR0TIbBoHPuYM94Mch438leRLEgGTSRgc9JNH5lO5gpIUkaRVgIyh2
GVc/FYhI9ZP/4oYogL7O4hpy4ft7pBfncmAXOg2NObKvyI0i6UUzJNetHRLelhXbz8lPg41If2Sb
1wEshU+s9bcr7qMUDlg=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
oFRFJPCQn61Z91okBks999ona3cAC1XzeoEwJREa6Y5vCOnNGKtr8cl7BGyxapXsQe9bielD3VaS
R8DuBzUWmHq9Ue7VVH+bU1BJ4mAfkah8Q26zrdvJjp4WKUJkWIBEczdySRbo+agwhKcj4UuS8Rlr
mCEkUM5atGrVL1aUEmbeETVMZvIJV3RRLeeWrQe1uPZaoBixmpWzwigfcMliT0M0G3lvSYV1h0Wv
RajKwrWU9zeWXMum9CjQQdZ3iApT5bJ8gEuwMfww3tqg3ZkxJ/siuWJy/hsIyqRMhlOtvzFGhEMX
q9Af+u8gJp9Fzn4YFceZYyMDs+qRLUehkgzlAw==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
li2JHyzf5QSszbS/GpRJxn/gUif/KhmzH8PNkQwkvztnOhKkFLun3OC67DAsoqlE3ygFUqCWAhmc
d3EozpmSYnBDBOt/SoyoMNUjiVgX21MfjAZ2fNwOQm5Qy77cgOGtGjQnzs6j4PQfuc9Ebn5rzsqm
lymk5yMEhSNqDXtxt1W5kj5/lvhxvpfGKo/bitEiApk25FbajjD0CaMuP26wJl8HRhQgVRDEUs4N
Pq+PXl5oHgAzAecRvlVI/gZJPRx5BfLgC+tC0tWQWhnCpYiYWRnC5Y3NSnD+1TJ6WTyVsCojV5/a
tG2OOWzNy1WbTr+i8EY3bo4K3jhtwhWQ7nREnw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XE5TTG6tMKNCGj9MuZUQemC+0MBapcCsaZ7dSNjqvTdgpeMsOeEf/IoI6vZFKtCO3ktny/T7mO4a
+JifPp0ojjFck+fXMQqeB831abzmtzYMZD2S6Aamtocd9rAKgcizHn1HmL4v4LdtputyAZLwFdLp
CcK16TtLdxhQOMG5HME=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
QnD6L1OxGlX72PPAJBR6ucjJokPNQH2eXfEsPgpJbOKKgcDEl6X+Zw8rRy/vx4ofleCC0vjgQVRZ
lShB7hqQnX4xmi+8O/CZ5gN8/D+SU5wDfQ/r2ia86vGCHq4X9lntbrPRLiWOhF7gFWpPEBX+t7LN
mkdEiOj2Rny9bEYvcORUjQrjXhKGqLo61LwW5WXLTl45h7xufa4gtReijrY7NiAUyYExJYLaEV8h
1kT/5eLfp1R7YyfpcGcRP6zq8/D7FC5qb2A11E4eW9F2k70RbWAb5cSqQ0TxH7NdVJVB69Mtr5j+
XiMB7LzGSYhc2csDfqV5Qpvj3O6uwGTq0NwgiQ==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35104)
`pragma protect data_block
PoHpMSVOjm6epHitWL2JU2kFeTUEamuwNHF5TtaVCfeA7uaCJ8xLWaCD8fhhbxWzThzwwwZPhG8v
iEzbUfuyjojSddPmhqLzMwyAR2+RpqlCE1jNSFEt9CBhNfRhBIXh4Cnewdiw/6o3tVU9VgbGX49m
xNZQi61GY9Fet3oi5gwgGDet65OTtZSGnktG5WZ+clNnqFPOIG0SRD6vsgtR/xu0udVfRjGt44qX
J6sM4KL4ITjUzCrHTjgtWnrbp65vvrHmgBXKseP8G5I+/l5ENlyUV2dQ2QViazGsbz7gEQFe+0Hk
a87a28XtUo4NeSJK/EOrRlwBQWvIaTB0cm5URn7AEyazlUAhVoQkNqh4sNaN8Crhg8jAFr844R0F
Npgy3xRDq2GjbjN4DY0Vun7vx22UTgOUqKdwX4yRgzaAiTk/DhAUiDxWuILsCsuG6NEWhiX/4D+M
AuhzwMQgTShO8PEzwz9CA66R0cA9uOy8utgMb/br2JkBGdetQiahR2Vn0MqkIXsxqXkTdIxis+JL
0CHizqcE3Q0J0BVCD9M4+oI4cV+F/WoelymfSl6L0Ldyl8EWkf8PmVG0FVeMAdwgv3d+BCF0hgX2
199VHyNV+qsL1rJDm72U0wVjnY3E8/m3l48C6Vv/rolAagh9clxjLgARggyvuCvwHn7Sh5lf2Oq/
4ZsDaZu2Wyrb/YQxi7Dl1sqhIZaMjOdmfPvwU23zqEZAkSiDpZ7pBU/2XUUu6ZZfTe/joZftFN+v
5RJXTKVp+I9cMyPswsyeUd3msEZljkUfTIQlDRW/iMAr/5EqL93eIcrokL+AdlFaynH0u+i6RcYR
m9JzSUALuAuwWZMFXQlYteabGTQo7n13TDYLtNd2HSkJLCxp9RDLKkIVrxVhDRBtSovrDQD0o3AA
EHTdnZApgplcYTJcPshMJi8pOGwS5rc39YezlcJgqHDVaZn3eZHTwFKaPX6ssvjSGdLEP+2gggHs
G7Bd+sJ/2vmsjuJ/MwC3uAVSQTpo8ILNMqGsZZ0jeHM2O1c7AtuUczQTEUWTTopi8mglPvaMVtEk
268FdxjBxirltaQPy4yid3mw8fnNhZR8OUrRHWP7SBsIe1bA/n1O/aGLZrXvl0mrYi0eFfkzX6H+
iWhuBGyc6FeqeQHr3ONCQ3nrnGHq3n8Sx3/x0OPaJWrSiwOwMp4KBY+rHhGh/rAefrTCqKB/7lcL
HK2FZCtUlxxMXoConlRadNSCjwvrtJqVRowzVdtZgqZOqmuhd3tyhQ3GphDeO392fVBMQFDA/RPv
51cewLpkmkQWUNIJSOW5Q60nCdiiikpav25H4DrRDYWG2OPBB/yXf36OwicMLl1DFFl3Mk0RzChz
eqW26hklt67cwa3gM8aU+h/fFiHeJcq/OufhDYVQncyBRkYyg1hw9cIjLHF10YvRK+X0SSDDJSAL
U7gWnsmYCDyKKh4DCJMDrJIOa6Na5TE0l5jwq8/NsWlb+Az43+JstXmR6Cgd/VCboio0IWFqEjSS
2YomXM5zIFmvSWAbv9COI+hccKsB7PBe37AFhAaEOt1+nQFQGyGf8JAlKNflJUcF1yfL/cYlssLy
RJs3A9NkCul7hqzeeYE4hg5Xnhpyb/KL57DjB71EI3GNr/GlWbhkpmiPigV9CSVfBEzg9FFunnBN
lUkd7jwrwfAKgDth//e+kdTW0xwbzjxkmcrB97aQ3jXgkOl5UF56Bdp4D4iKoJV0Omud4Qp1xped
tTk/SYBHeKFhmYYQKsNuuSiBYjj8xeIF4ld8l1k+9QPl+41t6VGgT9qn/hc0cRZig966RiefOXBw
fr88GXzkFc7IEYM1y25J004/zBW33gjIm2YdNwzBz146PaXl4mfCFQGElM7t3R3IUK92Njt3YlTg
+B/GRKDT3JgELRtpzXP3aQHztbvUPrs4PZvrmrP9ZlXoL906r+dOjEfAo3ZsV8HjcIkDjk47qm4i
jkR82dPFuAQz+e/D8shkWPCIgCIm/dhrT6JsSly2RfzK+QFYaz+sL78maJMDzcK4VEwMSByInNND
cuP6GnvbVHWELjc9g8TVSz5jyNaiCkCrB8K0JA76LvdFWpsSX6meYDmC64/mzjIQ+MZQB1w7i33t
poEEzp9eKZEtlDdzPUhZbeb/yh05TLYWHXRqJWMaK0eGj084RKOvf2VDSKlJeu90ijJ75TGJjwux
tjsCTqSgOR8S3rAfZ/LaLaTqGcRIHrAAbwJhgzEVurRq+SVCrwomJSV3P+MhGNyECRgyEla+NU6A
vdF9DiP8yelMGaXMDZ4j0fpvZnDX81lbAXHQ0lfk0zwWzXqlRlvFYgYbPFWtECtM2P+P/MxjHo9T
8+tmSG3Mao+gi+MnDys28s5T9w1MBFXb+nGFYa4PZKOSIus4PTiJZzBRyov3N9x87CarRYbs9ZfQ
fr+C83OT/WdQfVQ1YewGxwSxhLnSAec1BcUq0NkMbgKs4XZTtjTvWSPY4TnnGluEOSLrY8RQ2k7i
ljnsjfJxSzRs2gZyAdDZSZ/IpGqvdFUAOBZq/bW6Jelx5YvnQbqmN5tNiSdZ6NSPZMrCn/ZBmVoy
p/JhgyKpnim1BNMAjkJKVtYXDBWBm6zHn3LiPreTHPbIw6F/7qZ6pDovG0NRhvaG6Fh0GNlGZHfI
wgwjUZxbrmndswzyajJ63cTl4/DaNX6xsUgWtTX9EPy4+zDixVQKNo8Dm6VUbHCJrZ9bC33s69zx
BwAVTuoiC7a7nMMW06sStg0FTQKNtQ8GBGfs17E0qmzhykGT8+nmEdClKceuyMMpTS1IuXOuSLLz
HgyhleZF+uj9JWqzz+ybY61cFg8169k4npj+gVpmHlD5CnMkZq9uYSCSlkBA0JEAdqfgMRBa1Vbs
NVcr+Fr9e7hpziX5+n++TUaEhlrCedDMPIcW1z8BjRh++lPmkorXSCA9TC2hmuZolkLo82Y9Bl/a
InJV2ej081xVsQatjEEH2ds708BpJ6l/+4Ricy3EQ02T/2G6B96eNT9KCnRrzO1aYbU/79gFrwOp
FDkCKU257h10P6sVoCnqm9NQ0mfhAX2e4sfOFWiYBUZQRfVm3S3nU5fUQXT5/Tkeer2u2cv/Gxln
LjBYoy4BCSs94VxXKtr5A9PCFoiE8PBFv01iEuQDxaFDuaX2k9q1BwMk+k2CXX5uaY/ttwvnkqmO
m3qEEQyHU1dT1RKZzEMRfdadfkxHWdy0f2dQSOQ0wuQ8M6BYQUKKCLdWFz/la/zSEiGCVoxVTEra
xaHnXMO2CmVgOt2oR84WmZSRDm3eSqcdCb2PjKDiYswjLHGlOwFTZrBmwyGPKt8e5NRq01gCJHbi
W25P+tqbZlJQoBI0BDop/opb5PdomB9TVeKt/wcyftVrKoV6pPoNEMViOBvNBlsWpH4ip1zMA6ZJ
HO3bnynUvQLCe3b9kJdoRoKuMG1bt1odt2jrMr0lbWlhie8ol2CfJJltsKzc9lEp3VuGwAu7PHxF
bWk+80mJkE4nPlAsFluqY4nJ6pG2nGfD9fcl+NfPXDl6sX39a/XqzVmznGuKxh0GWjkf0b6JFyiY
iE0sj710UxRoOpcYISQkA8axYn3J4Z39uPEGi8vNJCBvrpbJGwDJYN8uovqd40lvWIOTV0FxJLmW
aN19tH+HWqUfpWzUY0xGCYoTkJdV/IzJVXOQM9CWZUXoUo/HXhT11APZ2RHQJCo81YRuE663O+lf
2PF1xKxos6+1cpt2QWAdt+OM2NUD/flNx6n6Gr3s83xoHmtQKDxDyQ7j5gyOb306nn4d1jIMQrcb
ox2T5HBpuU5/G7rDglwi/9MASSOiCTmHsROGwE5cJCFkX3Pe6mvmSR7cUdTEIgQE131WkQxcDFVY
UDz9GCbgmk5BaFu3mReQjl64hDLE0mRQa/J3XYnPWx1s6ZsSSQtYv0T+6uEKvzDn+lgwIjx/WKww
8oKlB6dPztZm/hbnxS4xVZk+GbHAKMXjURjtyFxw1jxM1ZofKlPdCDGpsQR28bggFM8Of4thx/6T
kButyEazQsArn8cJvmyrjqsqjNocUQUabpgBv3DfyajIjq6OM3Hi65u1tRgJUs6Ws5svVnGf2Pv3
9OvxRaCa8Ck2+JvyzHp7xbKjMmGLbA/MLD8q1zlzNDzE4EVHoSMSOWutDWMPvmAF6wITDO9i/UX6
0YiPQHVRT8pwSm13gdgfWDIJlK4mpyvx+A9bk8agoplsiC8zZt4MKxMUPMc1hHxSmD4POCn2GjSK
A0lM0kW1N1mto9KIestGDpWYNqqiPg/2F7p6bTOOKlhowjp10YyrUaq9DdeFKpwM/qQOpHbjoUqU
yxBCJllp3Fu+Ly129tWzbMxgc/FkXW91D26eI/ij55iorr/UQUYSZ0eXHSM5PM9SP2Zleh784ctL
VD6eK8yWQ6r3XUE5sq4+jP0leXRDQzNhOzQDjdQ2/djhmLeNgcBRyvlpbxp5P2pcGfDXHK+MZ31e
rzS1c/j2IzTxWNoaKVRXZIErwKvneiZs1hSP3q/3Zf0n2EBpVeoJAH7NoRyzVsrnNkJMeTTLEObg
NdDyFtDbQ7T24eYeJ9o/rou9OCbaMqvTquv5QyPqR/mSdnKwfgsqISmWBOoOuRY5gaAN3Fajd3/W
RP8lsTO73MApnxOI6XWvo3+eHcsEhoF3tIug37QiwM3C+t1lbHTSSXQ4zUAbzjRjE7Lb1oc7Ruda
z1YvUTYurnHKHn57qaZbt53ihrGB49827ekEAl+yX/GhS91B67ACSoOZLQ7KrxxmJzIPX6HtRevs
5rKLIJ+ZLXx+1B3uaBx/3Dhror+mnj5k/Bp7JmxfPwYafERadKXLZBxa8xo8CuSKilxYPbsmm5pH
IsNhhsGLJ19y0cLvL92NICwKNsbd3R0Hsecl/ncFudjqPAp4L7VjzRWGXUSqNqllj9DOROhR6k09
eRI10pVZ/UVQzHUETOYFpn2SbjUgLZaEXDsTueToyUaGvcWhs8IydILWV7MKRQZYrJFmhTjcCXNS
9bwZAHFLjBWLern4++hZ/GF/5R3QHcBPKPQETfXJVxB5FmdTcNSVCIToAnnbgndoLM2TO197mIMt
53DvCA/r3ItKrHdLxhBbGQDdVu3CyWKyoYsStIJxqWZ/wyx5vzupu9CH52pi5vPK1A7Y1pW0U1/f
nw1nMEkRzojeaLx7ashDrtK4WmGe2yPBiVVm2l9wHQiAoYgUd6/p2joXVAR40TXXmYLK6n873Ro3
wpGBUlLwQndNvKt1NQmV8wMKFPPknAAzB9ZYrQIQRIQwilVKXC+VFYq3quhxvukce4sb2gLiCjV/
GOYXgYjxhEgOWeMecDW/kTymTrbpnHi1Xnm12ZO0HwTbNNPofj7U6Z7PrAyMF9KEqKeT5I7vbWOB
tMTvXZ8gXcUzF8FROIyB9xKj5Nkfj+ZqE779G3DrvoAKdrFdOOURU+Lg9Dk7RxNY0Vw3RfEyvKQ9
PLB6WSM6LYOmZI4x/tpClauNkyklrUOcSPrsLedy/qo5cdkXSJAyRRRaw6j5kTUSoY1jC7dGaEuW
hAFlRciVFbNE5zgPMFHIGML98zrH2SAkpgw00+7aXyhXo4PXMe/fhNlf9gYl3tysA1fLts45kZyF
ENjuvbr6kPAqAybPqdN7EO8BtuExY1OWBeqI3XYNBTsowuAAvsL+f5iQ+baSgzJqvoWPITbOgRkr
oYCWmoyT/Wy2taaWrwTrqP7hzPsX6wga6lzk+BxgtzkeW/2YgMPyV9APX3Xk8/I4jVzuRCiVtvgd
YEcII2gCbsrnshInMlc3qOkIEGlSv1bGyfYZChxhnzZH9zh6rfLBrYb6DCDBoYemp6chlxMUotcg
ZgHEJbPcASu8CD+t1wbYvq0VDLeJ6TLhNVFWKel8W9Wz4YgNIRhdFVKn7vwxYpYXxDeMXvI2vQUx
xGUy9UDZKtAJJValTxV2oo55uJSIqoF/BgXE+Zs1EfCIOBvkk0Dyb0XwTtZU+i26mtwKmyCbjYfg
Y1Xr6JPfYwp92s7miUZrZTnL08Ekk6cjelPTkjpNR6LYas5G77MAOHgjB47a9E4quw2Bney9Yk9j
s5ysk5542qJnk9D2nPvmpOQLRNeYQ6NTFVLVP/Yf4cYIaEt4ejXU5JIGNGS95I+ECnGGTdba9deL
H06Z0YepIiGH0upoUxtO858jx+h6jbnXfvc45UClA4ODTYdUSpFiVoXRxbktFcjaejXIIzI0B/iv
neS6Tv1l78SWCEoE/Slk1BzMM32jOHm3efQS+q0Fk9OWHsjXQ5fSmg5/L4V0j8/RR7XpZC4bPXd5
gAmP2+81420RfxQU9NqyAkbQk9DTCFlym242sAk8/t6Vdgr+S3yDF80qRzuL1z8l+HKdnTZ66zA8
LnsFTOma1R5ciU2vHqoOZWxnD4U7LaDpRvAs963c0iSEAVdXdzHw3NWYZXNE9d3urWgLLkIkEVI0
BuwYNosR7LcK817nw+5ajhoFkAGd9JjRlWUq17Zplzia5eoYMFPAG70H7CTbiAdk41eJYO5imkR8
kBNosYoKXEA7dK+TJIxgEjpb2Qe/RDHLYfFj1FXzQBzBwcrIPD1CY1grtCs3JNIK0wfd+zU8zNUQ
o8nCWBBNOWWlk1P42HIKhLYSUJIiBfdr8v40Ivk+RRYH6vQ8Z578OjuC8IUMKmlG8NnBqWyfG+Uc
P6LmEkYFN2SgMxUidILi5sfevPUq0U3gETZYWtcxNYCj1vlsqQ12q4JThgAVtOfTf/WiLgjrrUHv
5N7sVEY31zmRmn2F2xmCJzmSzw1dYWoE0DP883Rq9c3hVtaGtpzT/R/nyxR3GoyRwyTP2Ub5FkiF
eKZYkQSZoP2bEpWvRbAvhw3xVChW+bhd112Jw0oXBiQtpN1JhIMdCmQQrYHuN8fcGzbeJBOZ7XYt
sqn7aFPk8EwY/B1kI4KFs7vEAC0HcoGrwE3pvreHcUl4t5yhXv/Yvyrj95Rzrpgl8VtwExp6p7eJ
g4a78Jdr/fpVo4w1p6YtFp+V8nENNuj/XX/btUTzhegX0gWqF62Lk/u1fMgnsZgao/T+Ag2WAHvN
KcCyORfNYz/AWjgKjus8G8MVh4wXMtCKTeaix8Hcp3c3akTcKDP3waRoPV7NuDd8P49LtGwqbwaZ
n9dFX+G8HIEycUmtNtNfweCn6wd7kPvKeJSX01r3GzwcSmzDpLdvOM1+wnNd+4GFR4IN26yYJEmN
OSMFru4KN8P6o8iUfn8vOXj+KVOvHhiDCCXzzebPHqKWhySvbCBlUtL/ojEUic0RQobtyA3beO1y
LiHx1nZ1vflZjyJW9hlzEcuC+XU65C40cvZpsqouou16KfAm3g92sWKEFhkNe9AnclpqWiiZdr0n
smknHMPPTbLxjCa/6jUjQ4PVGbb27C7XLrNVqUUcFBHmOm5RlyjzzbPM248XN/oj8IuhRXFxoeIt
GDwSWX5AaB3fRzd/BKhNa/zDIvuukbjKh5KCOb3K3PadcM/aVWPMlc9MptiNYMQ2S+BrQSrE6TgI
szkKbR+YzjSZ+xhxYMG3RM8ajY7g2uQI7MkT+JFH+HsrInlFwveep+/AueMet7ACic+KUWWL9px3
/L+z+LcX0/rScjq6WefSQANCfwtWUrK4ISjcaNsM50gSxRny437vAGZagHy2BbizJl84e4GOdjTb
Ljb9W6SexY9Nxe9ghqj04YAa+G1KGHJO+CXrX1DZWIDK9DSlDy7szD9gwFIADJ/zoWIHb2xo5OmX
FzfWoBRGmmcdPL5r8uLdlXU8dA0UWUXBtG6lQPa4UguLre0n6dPUeo65enEz9yNsHXBXyflGElgK
Csqxs5RHh2mIzJkBivspM27pZfZBochzl8KSclz5/HaNyQygDc4MQGHmd19pEXV/Jh03dyeOUwEM
lNk6FSd13SvHhLgbXZQgtJalhNj9JnBSei0W5zcZshLtjvNoZ8W4PsUXS/8WcNVfi/rg7If1htsM
9EdVFMer1vTdpU1LU0iL5KRO9jMw122u5wnas49QWT2epX2QY1ck9w92g6O8aHVyY1DzQ69sHH+O
j9mn7TZHE9ny0FUebh39C9FbbsJDdLKZp+Gvh52A4cL+AV5XvArDCjoQbYxdmzRaMm32tKW6SRaY
tzdh15YJDxH2vgGnsUZMG+X32vkt8yjIcbp8T7UneqpSbnFNBUTW+Xkcssn8WuBNfOxc6ybky7Kq
T8BFUxpvzC5mUEwPdcAMunzwWFmw/DM+GbmIyaTP9CjkO3uFReH5ksojbx/FPQ4hfOxeXt2s9goX
vTzW2+OcA7T4WBJ9/A2f8Z8pwGTpLZvTnMme4kA11M7MQWatAYh6rycuh6FaJedwERXOC6aIqbk+
FVoyVot2FeebApgKoe52MIhGJr2mSZ4amRRCQUDh7CaAtWicof/5lwGKH5P0S5l+Gd7K63Gy6TdW
U9e/RYqFBuX7y/Dwnuwe3KoYKaJOY5O5Kt1ZPrDyo0x8UGj3UcFrCTEt6ajeFtEQYsb3NihH/AHv
CI4bob3OqLxuaXlKHNE/GcAxTDpjE2fRCvm6VqqOq7ETrtQxUyohf73z8N9Hk0jS52PLUbqiFj4N
/XmdxRa/5WCmujWaefKDhqSh2VrqfQrwSNf0O0S3pOksOTQOoTuTWNuHYO8JW+BSZG4KqqHSDLRs
D2lb3xJm6ArQi3pjn3mFCYBFmDU/PDg6Oh1V5UKmfPISeMtz/6L++zTftDe+ZV45v6vmMqHTrnuS
iFWKMTKkPSXaUGSw2QyDgeyc4bvSgET4tNEb/ffdJ5CGboSD1vf2KHgpi5soQEnT7uYr1rJhFb4L
emKQHsUBsZRqVl6qeb18uwSs8TtI0QNj0NmEVtQ/UCasy1/i1Hb1KDRhsx6Qkg2QC8IfFqULlmPN
o3RiQn0EMQTwTeestRgqDjCD2DdEEjAPgOul2eHfWBrsRV2NKRDO7JS8llbqBHRbEaIW7b/SS+lv
cvgtF986V1u/FdBkvuqbnMd0/iwKYlHO5IoWsysD6rxY8bASmOLDLeVFYI21hSvfvTa+ZnG7D9eL
jJwU5CfCLQnEwee2JXMv+PqiNVz913u4isPfnNqX6eY/9WTVjsZjpdngIqcMX6IdpGUTh3kfKqM4
IdPkmQIHhkNCRerSYTncgtF8LVHxnU1o39LvBc1YKCqe6ciT/dWIxZEkVJKLN4jXIkewpX5Vzs6O
YpUGudczNjjcFqex9k29uDk7ZKteSkny50WXt/IFCbKD1equZUXNtsNRnAXizjNJM8ECJU+beTnk
tTUZRYqnR3p3HwgNJUqUERWYTpKakRG2ZiuHM1zlSebCRK9CEvqfVBn7vqLlFDUmbDVh7D3Feoic
kYlLDI7is867it6NzgMgufVr1T8vpxG5LrzYRJ0WPFTcptEyHUc30HFhrxfmjZZGy3cU5iumD/wa
0ICYQMQfXis8av0EctnE9KlxyOlE65U2Ztsjp+3c7Nk6apaUQCtAX7L3QirpXvo7aZCmSaAcL/nk
uHmeajesg7uGLe2OgXvTdFoLAaglUgE7xmTFhJj7IO+Ou6Uga1vakDiboTQhySGSs7xkI23hev1U
P8Q6YkpMud+gFl2nVXOUtY/r2WlWIlCnKq6wge8VRA6dDEGgRWumh5GgYDoW7MHmhyFuc5z8sFWs
muKauIVbdpC8x/wyBLZSvWapxYUQovV9+h0sFt503us08mZgmHyMCfUugYlnjhnQWXiYtLTZMYd0
YjPCagNIW84vXpX1rnbeHmAPhx9GWNV8ymqulGJJuNA4a6HuyfygzY8oxlAOk0j4dQ68meuLcgD0
bHY56DnlwkDZBK11NIEPOOcnXyX0WrWioN/QolENIW1lz3cRvv/jGXtKs5L6/W/9MEyIQzwQvTDl
WCsKLpPMg7xZouREZAd5MBgmtKp9pl2me5MHd9mVYOEP0meZIKmaa8CCdDCyvVaZJehvM4y6Wz99
bvGW3vZQwM8TNdZzpzlW3Vb9JR3Q0KqNpXuotBNAl0jSk9e4VSwnFzRmwq152qr5FSB6S6TJcgTS
tXSCBFX3Rhp+ptbgcUGfCbvljs/eQ4DhxvgewCT8jo1i8hbOdnd+onXGyzt1fnqLjGn5IqRDsYtj
Xn9jo1NudV+OLTaPvUmtqyQqMhBmE2hFyfv2m6sWe5G4O+xjuGF3W41xbU0XBu5Kf4xQjpsFLfmj
Gqg6AVrjZNdGHUy0Hbb0dW+E4v+pXnmTRml8SOrb56nUNSClyKjW1mdRdTDrtetnwqdDCe7DDheJ
x1RR9cjvcEiMrCJpHg+7ZdEnnbFhpDzhzEZZD17tHuBleP/ehQ9bHQi7c1nIwkDLHmHyKOz10OUj
FIC9dn9s5yIa7eesgfTEmfjRRD3vcvGUMFBjH032oz8lVA9EtxL4RaOJtQJ76joI6w8+JtBU+zHy
kFw1rvAPkl/rApbkgf2hAmrxQKscbH0awzllfpVsx9+PaQgaIPMzl8whK37hwP5S0skODVN0Atqc
fKzoj/1t6ZJox7ZvCcjaf4Fq1FMJPzp13B5oJfz4eC8WfcW9LPjHQyEiyu4JmcAsEm9CMZc4wmLw
ONIHcb2n0k4+G5EtJ28e25oQ8+HmzP4JydykYz/8VAAOxm7aywPJuuYgQUjVJkdgnsf9xV0W7oEm
mKBUMAXuuRVcj3Wo6+vLqCqoQojcwYBO3gwp9KAI/pwPjjGU59yMQXPCMFEIqKczaP3oj8sojYZw
ErhIFr4dCY3vcgLRK+yReiwT+uyMKbk84e79GiOZpZ3+tyulEnM1XHr6dOBkCb6o81BUwgf8T+VM
80QYJfZh2LHzsQ8aiuxJXjqw9WVeVxEZqjLDMSOA1rZ2S2pen8sOP2vEoHWXtTm/H4rXwodqDxcx
1+zos2atO8qJh12gHoLA4LAoZYoE45LnJooub8y/e4R57SGlVuz/OdaEO9+XTkjp74EXIyp+j+Bk
HWtMv1+70siZM1W7FXY1Dzss8qYkF44qVd9T3ITj9zETflVgz1NsO4oOICpExOH4oA7Q6ynNkUpu
EtP0B16fOS/trXvcKZ7zLPecK8mOCk4kHMGLUDRBSH5yBYR9mAvMVP+bH/SYdDkzfB9EWPNRk3t8
A/y0r69+f0PgbAMwa93ONis5hYhcMKvg/llP7KkUWSdDjK4fLfQPc/txvyQ02k4B3TVWXjQ+cKAM
Nxq3xiY5LAxSCJK9p4DC4dCGIxnVqt+js9K07vCfN127aV5wezr+14kI8AmI5ADoSPMQIMgJ2liT
ulG3BvBLVeCdF7RXW4mq2qJtMVQJPnUzLLJuFMVWJy86sZISyxFP8xIOP0wowoptIP9Zdkm7kWKg
8DgB2AuGC98z+7WXLV8TV/rzg6eDxlItc8QLP7cpoYkw+CoEwcJNOWKYNhZzehu79noDoZ5D7GEu
QyJg/3JS3A7Z6mi5wdpWVAjJyV2J7NK2UZzvdMnC39NbA8WlVRwy7OiZewHeQLNpiRzQtZsFEVrw
R/fQpAYpl9Ig9fOMLzp+zuB5Bu1erLX4WV50N8gNu+BVNVXJhGvWZw0VVVTDTXQOXQu4Hg6yDg93
Whr6jTUly75Gz9aXsTD9R9e9tWTINrfb9zzH9SjA68UcAbsETpwk79p/UpMmGHt2m0eHxlJVHcaq
Lv5RAJHI3fkMgf12Wq1xZ8QiHnFoCnL7ltDqvsa66IhvwfyirH1V+gPtrVE0jKgMWLl9gaWseqB8
0icn8k7sgQIdAU5yGVK56w3TTbxIXvqqKbcJbPYFxqIOKMQvAwj70Yf/ydVSU5OVpfqugucxxZe7
bTU5tcz5CR0O6SK9gXTyMChbA09rWGYkA2Oqu5jv8Q6v3hvwpkJZ8El2IgI+VDFn98E/2Bv3kM/z
VwIC1A8T5gHTsSd7HPCxsgRbcGrFIVcHKM+b3MezKnMkCMX1l3EgYUYb1Z1yaCE8bJDXuiIj+K9E
J11CunZn1LT1s3EJ7lknz7K1cKP9nmE/ywaiuvpGh8dvwkqqlw7jDCf1cBu47IbWg2LOizzjvSVO
64kcE53qS8n8I5vSqc9+z8qVwj3ed3BG46Ktmi5NCcP034vvF/ldViMPBsyt9O9yHH2m5uKqu0os
NSG766LqBXC4R3B7aQW8J21SFx5MYeLyMRnrywoB4fm4t6elcvBgLbAtxqjhzWc5D/yO1WADLPql
NZVcwr3LfTUdG7mZ88qTiUETiPObxGxf+Pl3nW5HaXQT0OEM1QXAUSXVYy/6ix+TamHeMsEY18Hf
e/xFgMJE8WccAdxOD8Oa0Yk6cXeaGmih4oIsQdKfzFSsrwk1eX23XAujKD2sK8YT5hWo1hXGVYDz
FX5+n2Uqw9l/UM0kUcE/GAh3fVYnTAp1k8oLV1OLPtUd/J5omJj8/tqMcOq3yxX7xa62IeysVFoh
9+kQLaKjjubM92kb4/fqrngYQIie95LN6vzJJTCqvpD8nGX9TC4qx7P/4IWLLAC3iKq683PgZWfs
dFDqaVIi//rcl05QAgs281+qJpdl2gi4Xivdr8Ex0P5xskjrkH9HIfr/yp3nxuT/K/UY4rMDcYe5
Gf/pJvUE9QTid4w5r+1zkc5WR3Fo+7twP3GHv2sg2Cxb5tDPhW0pvnxrxRumpRy8p/592RpwC84w
YpJjQwYQkPgimLYux3hC6CwhC9/7+F0vp2VLNcxGICqDk1o3wAMMkqrnb+AG0IKqhDX7cxjYmJBd
T9gBTikK33A3rB3jWYal16Jc4frTCHXaNn1MO4jug30jGIQyASxZH96SzPWSSJuph0y/cLulyaQq
5e6c3378V7E8cotGdp5SyPBHH+cdgFrtBE2SA9WuE0JW3Yh8vXxZgOtItTUr9povhS+92WJQjRlX
tBsR6VsfK6nmai5AT08HqbsELoddpc2ETlDvc+ISygtUyGI6JsASkK5+bUG/Hn4kffgys4jFHx7j
gxAAci8aJCmNpR1ygVLZ/+99rum4QDxOYoyiwOSQBfJeqM1fvIIy1MP9ryWp09dgPHT0tarFafan
UFuoKJ/QmzAdkFpdY0BmD7yREWO5HXB+Rnn6X417pmC7kMAjqDWiv2dlVa4+d6qcU3Y11h2VChGd
KMw/78AT1W6xQUcJnV9lWo3F/mffklrjF7aXoHS6R2Iy2rJpMO5Ua5JvdE6Fo32JlnflKWRDOYfU
AvOq/DMZ1J4gudnz/0N/EG4iL5vuL5SAKco0xiegDZKmP+n4hQkOnoLjkS6kpvQ57av/CBemx48H
QcJcEwI0/tgzmrX9dRkk7/+wvZMqxDLySXjtewRA9c52BPHcag2sI6RwGnrdVZir9sz8hv3PL5eU
b5YleFRXBaYLFAL+TOaHtqHy3QoDTM7URZvr+tNnH8VmyrG6VSDpr2ZBijT8qcZofYej2bSa353K
1rZ3C8GpT+ena4nA0pwkJ7uHTw9foidFNGNsKci6gcoKftp9D/Yqh46yGuUAJ9WIuskamUqJFeGm
ce1I2goRqRWzS+qaOUjGMLN8wDdK7e22kzi8gDHcdtPruxJ4aL1aj7UAR70/7swDNK9rMfWfhfim
L/bdLpJ6prmPjFINFbkX8xW+bX7FBpi46y8C5qR0F7Vouk1pXXKVzFFAyydl06e2FUrG7vmAtx0V
zwrRiSg1xjtHjCfyu7SfOut66pVCWyi1+jQNZ/5cvpig3i/dh0ePfcVbq3+Vu90vKg3gwuz2bZAB
03oZTpFpuRS+LzBwm3wHW4zLcuz54iEr0TJfczbp9oXYc+9HDzaN1RINZiecLfG0tfqhAe5pC5Vy
XKQ1dcHLbzw409YB7qgjIE+gAlRbil2mqjgd3dgFmpz8Aoyo2LvGh3F2BZ6a8UKjzvJ54iRsnaSL
mR6bjmbNdDWNROFihXzuzSglPDqNSQTzx/4r1sa+3Z8zgDuiQadXJzH4URM5EU+j2kTqF7BvbWjx
MSjQ7dvcAjvEeOZBeQF6mG2i9XpVJGCt+qKjEuehPuVXR6RXjZPspM+K6elaaAaA3NeYCuX1HMO7
UpoRIvZhq1sXSS586WkEDqKEIxqqW8X+YYGGXmSvOjFEjWPA9McWxWrXk3vpqvHRVzaoV8V+eOhL
toUtq6EY5PDYZ5qVI2B+FWxgewmyK/Gx7iV4wOqfZGuHJ0XinfWzFva3A6dSPjvpv4NY+RcQr/+S
v9enJu+qMqNdksCxeA/A4d/sQYfuhKhWmDeetFC1oFBUjIsLEQPm/6X2cf/quG9hZ8YZ9mR6AarN
FB4Kk8LsK3YagTdcWbp2Na+bmDC5G2VmqzYjtsXBR8OtaHFD+Bn5FQEhrBAt3X2H+ENQanFEE36R
9ekcPHB8sYD6uHk+JUN5pKYZKjpfod15shxvYTCkPc87Tc59W34TwSMsWrlfuHLKZJdkTf/y5U/O
mVoZt3vFheQ4QnCesrEhgoqlOErPV3pVTLEyclDXJYcwRvfPYwPP7qUglnbSv14XetE7cS1phwRN
bTXiRCxEINurYf/mO2FvR8FyA90wye4DHF4A+F5Qf+SsrronidFObGxQ4SA1AKuElYMfnxfgbMr9
N7rGpGojy5zCFCibHtmY7KFx8nACaiHWvCm/6hr4l4eJ+NqB/PbVzs8FGxWcJTprLrm/PFoNLEfK
hJniw3dXx8df47KL8/lfkWUelL3S0EE58xrQAx2q6ycewurHGH4e5wt218X4VTFIe0aBmpLuAr5n
+ALccpGGSQVr4RqQOFJFvPCJvlAtkZ7vH7TNt1M9K6798dFH1wMQmIexeMicUEFvC2F/zhzTNATO
qPhyZN8Fjc8Eza/C4ofY99ZtOqfoU631MgrikOhLrTZ7BXeMQaB9Rbj1WVT/xVLPXFBKF6e4PMAJ
h5boAM5ABWJCFagdzXjqZhuoOCCKE9RNh8GHw9O6OUb+h6YlvOKyIUMAEqFGI7v3stSdm2jWV4mS
8dx9U2zmMrfURfKQhzpW3Ju2+F9VPZUqR0etx8swefCbHnqOtu+/6MHegJjEk5zL6+rYnDlZfV/8
/GcSALi7vJNUOSxXAwrl93By5mw5l0XtiW2+D+9jYqlDqQ0AbYbUUi+5aNtJQVp5mnfdURJmEIkJ
GLUR4CXpZCbQ+4VVAhmFB4n7vuE5LW2BLLta0xdB1Yav2h+PdnlZ0Xmv2okC4U1TLdLNN4hsGIxE
QFh6Ih7OcfcxKXB+lCErYXavINIvPQcbHTF4s5930G2di4iKGJMdxo4Lk7MWB69+hTRziYcA/K4n
A9I4czcFCCHF49A6yr35+sF+UPSxnw2G4NH2JY3h69VXc/nxAnCGoVukrr6Cb26KgQjPPygep97v
m92lTk2bcC+rXCJCWWik1gWqWJfsIVDQKHZL8EVxRHOO0L6djEE6dGv3Xbt4cEdLeQDa5XaGkgmq
g9g/8UVK1Zjxs0Pf0lhiLIh7fNq8P7/Mfe88d/Wdqma4Z6oLaUx5egbTVEUMk/6FFOQbliAoASIX
LH/38TurvOLO+RFjzOTUZhZLSpfdOHK6g4dAf+pN1pbD7DbioX8IBf5E9N0dUdRzGNn5okYE+i3Z
bZpg8ILdQl7v+F0RKCu5XOg32/njLCWnpxtSQE8OCDUgymx0IDCmydfXQka5wFHTWnhX73D789Np
eO75bPVjYAzcK3J7O/AQc8jVO0csTlp9yXxMrKo3Ln7V+8XgdCD69WGYo6SdVj4jS58dUgo8A0w/
MCMBTOaoOLoznYnMqp9xvb2gEal/eECxTk9+Jcj03THp4pOvnRYn1BxYMM2WVOq2zI2jOWNV/Fbx
GApAS/rN0kWQ2mjhHI9Fs9KhZypuQWn+SEFX7Cbwo3MM7Irld7rOIQ8/C1zqOGtOm9JvnCBnVDod
+RCm4vpbD0CevoypvF86Q9RAKsqH/gD9PwoZLZyDBi2oJLDpyoctxS0CMFLeJFtoYNH8Pyk5UkTp
DSAcstO9tdMRk28snfGd4VBo5yRZWNjM3IkPuSgeM2XrrLDE+KuiqZYtGCTK298SNKOXc+08z49P
leNa/NKKXu6geQASylMqSEO7i/FDB3DPGHMi3sMFYjVYTfL7t0mG5nX0eRZBaBzJTJhdMRwDWX2Q
gDTiubiHPhChI3ZxDRsba4C8JjLT/noVOxpdklqj6K/95sSwRz09Br0MHfKfmacc6Tmudd7Q36Gm
9XjsU1whpJK0zJ/npjg6b30wAumpIEn9vy7vXHWYw+7sZ0oa3NkarrIBaeSk4Jsy6IXRBdiDtZCA
Bv6wpSgQXASDoMVkpfvibJP02N0ezZbglz22ZoUYP0hV/u0cHuqkjfLFto0RlGt1i2ihi70pTsr+
FBAX7nM6/PhUJo7neExAUhw6/UxSuRL+2Z0AQCAN9zJmXzlXEu9gXiCdohplkxhQdY90L51GO/ws
Sj6xqUTzJJ30BDXaa1Bt1w7ZVJEbN/bkmpXSnKpUhOqCRQBwlDrRMYOPnAe3CHYCm7/ydYborL/7
tdh6SNWdV8IMLbjZ5oCv+dyGZ6q7hnFKJurtKnr0H5pbTg6g3Ll4u09B8a8cAluzByABwCAYWylp
p34fuKfeY1tItvAY/OfHMe1QH1Zb7ucy8MbEx+IjRd1Fgy22ced/Xhz6me418z1FuIj5Bodj3YkE
jXKL+uOjbiOWwlWwnH34Tz2MJ4dA0UvHZK3KFmlKsxSIhp3ubJjlwd3dC9RbTMrmnzZ0mepc2uoK
MMtRtP/iFbIjd56GU1AFuK0Y544lxVgkV59wT3twjFbvjXum5fpehqaTQoWV+rSUMmO6TzpqNDaX
8Gx8chybazB5xdNoTqVk/soSkO6x1tVsTODK982c8bsGaEAzRjcr4qidzw+kzQd7sLGFwF5UHoYU
rgpNMAm46e7aAWipcrhn4X5xXZtvCHtnAnsmiZ9q//7gYCTbSU/ZRyz727EU4wVUV6kTT7T98QU9
VM100uqgaBKlsNPkO5BxmG71BGVAuKqPRaQuHKgA05nl2+Tg9Q1yQbEIaHGCivz/iYaYuaW4ze1u
QDdcegliK9ZE0c31L5CgMl6F6Gm9CSOTzlUI2S3Oy/ErsJh8v3tf6r8rUfpVph2NtrsSHE4yRKeR
YUGv+B7zxGUw89bLUx0KzAAe4TTG5HDcWPzhU17/HwJSUmeyN8mHNlFWehSaidOIIC2WAs1BHQdV
h+1DCHwWf8uYBs+koPkwy7UEve2cPf39LaCLIeXsCU9pTMGTLg/ac7eCZ29fwTblSok8/d4GlnHH
frcdzxUoxpWIVfkDEHcL8FDThDgynqbO7NvOcCARpeTpaV4JSaJngeg/OGNmpsAwWjUXRpzxLKNB
txrU8OY4UrbXVkNRHUcA0GXS4Se7narYTiIhCT9OGu4TeeqhKe6sIfaoulC787TXgtE9g/OVt2qd
U4aplgMVTnCLmQ1FPmvt1pcCpK170Zt+ximHQgzMfiEgH+5tf3Tq9f/J2EWnecZVRFKWPZjZbI3/
jpnTJkKAIKlN5M+T6ohXFlEd5i3f3lnjJZzI0XJfijOa39EmiB8i/YDDJCASCqv5tyzl+39BFOuB
tHAAAeTfqq1ThluwFZS7bSB1+heMcJKJReXjhgmEdqEwGROMgl2Wu4o8m2liYeIHBQ7F9baYemJx
srup2i+luFA5jlBSh0PSGKZNreZgU4jYnefGZqlf4aiDvXfAt0yXUonFwQzdDwQtVzpXc1VscREv
aiIUMTO/GZE760lSCzgoCMV3zV9+28DyGY52wGk9BmUtCQagCdLkmrnmvGd7kmjjnJM0IdRhPMhd
4U1cX/pXaVr/GCa9gkbCzpoNTxjMoBL9T1AMPoIUeqjCRrv82vR1PCRKEBCBBPRr2GAlIdmZALIb
qC7lZROmyTmHWrPYHy/iSEvtvxv4/xf83B1YhJ6Aj/3FfNeEJIWkZ5fThZC/C6sE+RG5G3ouKj9w
gYu7c4F9Gs1hdKpsr7uJqDhBfsZmBJlOAWowJpYCOP1TBe3V+nJt9eV97XDGT4tRp2/U2Ic4MWz8
iNlOWS/EFvqr6FWFo78yTt9eSjONVlw2E+E/KydCSMVnd0Kx4euJhkt4Dx9/syol70F/2NTXfopj
vtWffzQzgmHqE3Zz8MQQ5+0Vkr4/EDKpHVXJ0C0S5Sn1ZAlYKBkGdBRUc9+1CPcyGHlHtmp2jByc
W1SuOx/D/EP/0xRy6XEwhLwEgD/3oBlsaQWlJe2ogFXDFgsp0aA4OX1bR6FTEYsCNCHnSIKicVm8
1e26vQcEd6BdmuQjpgqHAdXG860Ckbe3T2oc3ZSkOwqd2SwzICb1SGXxVQdeErYg/MFh2v7gsgLl
N8T7GdX7DoqlHWXzoVWkEusiz+RLwnCQQes4dEjuHGz6Vvg+7XaJnK4LhkqFXysmH05vbGixittG
e07zKWToe8ea2mkg+70Dl0R+hlXRNkrDF1XZpFryuRV5wPqHhGTib6GeQTkujh2jkL6Z2AAOi8zh
Rv8fh7w6wnc4JEwOg+SgH/qkGNwcSRdb94JcfbsquW3sMh+iifAIsncIqgOAx3v1DHKG+2a+ABHn
80HevWfGyjo6w8YVWmMVW/4Iw5b1XfGZqz43BjLYsxyID8mIlIHOIBGCw5bMOhz7IuQpm0CP8KED
ERDIrkpph0bGc/yVZyzNpuIcMD3idEA3pQv9BJz3fwntZZrggl9mcLgL6EFB5hf6Qf04J2tHR+ci
fTAUaHqazBoVr2QOyQ7mnKaeWqOMSpEdCUVRnTYJoGGTj3KHk4Yo5Q+McJcWBSHo67bz3VU/KM7q
8SEp1VR0KSiLymQF9EjJCKqKHeBmLtx8k2+nmo2mMCnjOYcScKaTmLG0zKX1dBu5XtBiBm3F05pV
DJe9tz3TW4PgL6Gel7AVzC00M3ucuX/OMGlpfiYVpqfmu0L4rqrZztnOBhadjIo3b6veN4Vi7eRr
TFLR3yMaCz0RXAUZt9kfDdiKXBYoN0S+T3RbpdyFv4FzXb2xEbF5En81qyD718PGu+12HlGYiAj+
N+G1EMJs6VgwLkC9a47LLar/qTLVZi1kNUDV5qLW8NzQrsI6hIOVaBKbWNViyzBrJQHPIKcaB25R
ea3FkUz3nLy9CNtuNxf359RkDNXZX4Vvd+B64272Yo/p6fmNKo8QQzXgY2WC86xjeA3P8X7G2Ly8
pmihF5mt2GQxUc4D6QM7vQ2xD9qHQX48w4k3F9y5sAVR72T7A5k7riQEKKJoDkS539tVWivKoGoG
EQGGSO9K4I5iBgOkZ3yD+/iFMSS8hITS66P7icX4D7dMkyCTRh7slii3lr86qlaO+DDQaxts4Xt9
3mRWa6CnU8j9A2a1PoF2eDKI+M+tVtyw9BlaJYy+qJJiMk4zZMzJUBrKzmUJJZogBRLO+gKUJHJe
+6nr3UbVtNf/64hbbdYwKKAprDYiUnV1pRhF519qg14goNurHcHONlUCqfkHDIpptM7YpYArt4h+
vQh4GNXG1AbKt+2gUBNd4vpUvSZ5eO5Kcet9P/aJcIzqMZr+TVhZuBQJjR569fTbCAzKJ0QVveY7
mfrhvXBsXcNg1O0V6I1E+UdjC2/3f5thnLQMoYP5dPRvw7cDKbP9PPqgOPP/RbmJin7/OXOAklaU
YLa3ZdIyBNW12uYrKC7zPXYY+j0PijueN9ELwCe1CGseiCbFL135SCnhY2lIlquLb6jnR+qDN8x6
aUc6qXJf/qncGJe3LEYW40lcMDdeBRr+8tdTqsB+yD8auTDAp4myebwA/nu6Q2jsoHXySNy5MVd1
oHxtSSZ3fZe0aG2k1ywaVVbrdHLOrOSzTwYw24XDlgBLGn2wH1c2UiEOEYCALsWnFB/ezs89s6QV
Yeq+gkB+QQ1ktzEq7CFQe3mdpmHvWpjq1Ezg8yv6eG5dPpyzzYMzz6EhgThHrd14Jo5wt0ip4FeA
SEHs+kqnSdmD60j4/kxgo/viX7zbe7DCpa3dbZzKq+jNH5UsissIqBSRP5O1ooPbQm/LRg8D64zy
6wmGP7QTsLFuuGlJJS7MdOJcV69GjiNpc4E7LlPaN5Ry4vLykqrje5puI+k079PyhvBhim4+5vx7
w/hvza0UDYISSMitp3PTv9tfuyUX5F8HjK+6fa6izaOcIrjdgsPp5zXuyaQQY5zz6L9LIKWNHO77
FbLqqcKL3mCnbXOnfRWn7itHBHNjkxjwxIA9OS1m892vpLn8leh4u//IKQgTk5+z+wit9Z7okMtN
Zmx2BIHte2Cig38hVBho4FJIqVF5W1XV2ZQTnLcFJjjugoiVoVLeEZWqIqLLYySg8OIyD2FthSlM
G+ag5505+is3gJkOh2JTLk0udiaXWxEuoCXoSgDY/sCpOd8qXbwrwP6/u4sIPU+rukXLJtsUL6pw
iRQx076OJVhRWkPjjaYTT3CBpZ5di85kv+jMGemMJFdC8uAD//NVO5HMQysnwJFjs66+wQ6Q0gwg
2t1dBf9qRAT/uBaryZ7Re5EW9miAQqopYri/p9AjTKB7BXzdbGD1N4++eopjfZsJ6wZ6hoTcga9Y
qcg1gzITGXqYMMarW4jzIJIUgiG7CLF10DQN0Z00ZsU2SqIa9Wqr0ToEUKJ1OAVPXFw7TmvxLRXa
fnz+h05g3GnXJ9LvvtpL38e454keJq5GBhslbGdMnHTQU4pV02r88rl+wEbYvbbm1uWPZ13NBKpq
WHSS5TJkeHCBHuf+iPKEYE9Yk92rlz7vl4acMMhHm13P4mGpfVC/BOSvOMozP3u43neGHwXJ0I6/
ujJYFpMCVcE+2ZmNp59stwwYUz/EC3xRgKqXKBo3g9Esm1rfuLSmMpXa0f0gC9g+xi4yokfcSKDN
lyQnRuOjP4fzH2mcbIdDcg5D/WAyl1r+DNkT6sNBDFlyaA0Mh4lAjg8ibm1b5zU+JVXwIoBuvftX
tQmWObdgXwlxhzYE0P2LYz2P0hc7HtPP1UWa+U3RydeIf7wRgGY9k796tFv1BSkvaUgui/qXpjb5
2jlndRRlydmhB+/Z6yALg8586S4nqhXXRPzED0dn270zcxkAeSbp+ZDGoMv9zuWltTB/tRzL3ZQ5
oY22SB949I02WM4C/QXqEAconzWYJXOocdJ3AYQdDxV4McThgBhCnVZ++b5KUyYeFgiXU9Ao3rrC
fpzQrwpSZidNjr/O+tO8D8uRzpZKKcISWU6O1QxQo/zxIrw+R8dB4DuekMsrJjxKx2nU7WCm+xwB
ohD2WtSEl7umX6pPKM+2JjqbhOEy0yLtCNmj5NX0sO+y4gOSJnBLmxLCYZq7UxxhFi+Bu72ssCG2
CZe/6aqoxW7DvJ/AUK52Xj5N+Q0JrpYXto5D3wELluC2LBVIQ5g851eoxY8nYP21YCLcGM2pRbu6
UL1ECRL8nYlBKWlF11057vO7KkYSovljL6R4lTixr8vS50kYlh/RGJE7djj3DkloLqGUPgub8zwe
Po6t5Tkk0z1sAQ9JGYZ+wTE8Fthrgr6x35HPckXKpGLLN5P1d9VhtBxvzH/5jBeVyutzWNyAaamL
TjZ+eS/68TJF4t7yPwRlT/ciX6cyrNuNdwJts8Q5Somvt1oaFTfamzOsc5/gsQB6I1UzrH0wg323
aVbWcVGwGptzaMkQ/XmerrtdKAV47/yFbC1xeav4klyLEvja4crimU+by+BJ/e/zflkgWLXgmcAy
w/aJByjOmfXYMdSJUXN6jictZH8Cy8tvrgJs8+8plidbWZ9mF1wRF9YygXQ2ZM3HZqP5tOg1bTxs
HCyfGIdl9WTGS5VAxtMN1CyQxxIjJ6JT8hgwinYvp5AAZP3mnf3Oi36xvznKyCX28GrQCVjuJpAw
jXHy/wdRTWoquy/GwHv1XEIVTquZSX+kBNZPWv/ETptOBN8rskehQLXD0PKP+l1HMoS81emq1QG1
TSJI240wpZjDP3Xul76tJOeXjG+6C/MwaRfkaRTLcgaUec/CEodad+mkB5DlK54yjSuV5ehcPbiY
jMQDaMBVhkCHFNGaD6dAIppy2kp6BV4M/fyUyInJRDgoOTM5JjUom1sxQcJu38qkrPPwOvyS8lr5
KDCso0lqLP2StwEDa4oKxPbYNYRvccvDMjubNBPIgq1StTeb+CwG+T+FBlmV0squ+CTQ32UGiLKI
VSIqkdOnLbYaPI139vLIPVTCTcEby45dZxQnOFM+CEGOcrpWqmmdCb9DFZ/tY60Jl0y+NZ1PhVIV
MEFnO++oSnUK47GA6NkWQ+E+3gx7T0lR4TdcqHjxDnDeZ4RdVPMx/eWQ9dfKQywfBJeN3jEr7tlq
2RaupdJtLiQsZtcPhpCpXZy77XEQ6tHpnAtlzTq8JZg35JGIiWRIYYyldlc6nbX87ZsjDCF/5YCW
BRqef2jVZfBSlLcm3cY6tCHZ9oigU6uihb/6BfFbrN19TtRK0Mtev2WGyhRkIYg/oyUXFBFJO3tE
z+IxKdzwPVgJOt4V/3/Q4MvWeP6YYn/95ji/t1HxhvLyaNWxq1SN/9TgI5U++5XhYcw/iY1TUZTz
Emm5X4xVC/f503y7RFgHfSvZM11snkC5N3Oolti0w/pWYIDfKHpPYJymVmYnr2VPE0WKndiCXdYF
ZDXwZdETGTwgDyxw1NqDsXhkFlLpazMUB7T4kln9uxukIUDvn7748GnDENedahr3zTRLzkQYCURM
CbGAU5pKpnQs9I6Y02g1gu5cgnDV6+UpMSIxFPkbYn1amBQyPSolsP/Rq4eIdTvNJyo9/lWvPf98
bhWNOF7zELSMXa6CppseN4Wny1zUMcJO2zNIXL3uFvpY6kKUfkyKs5r767gQgh6DE/uJki+Qt7wW
jZkYW1dQNyLxtjOmMNRlD8px4rPexzsvNXFtoy/ViT1xvDbV7kgyeSxrnqEEimIArM4C/lybDYcZ
omuP8BTb2dChOfftZGUictLy8zDEwf8hftT9g77c16BPfQG6UtHsDQKJzM0Hv3Qs6Nq7pxPO1BUW
XKnh73W8MnuYI8U8BOBVOe31Zwl6PyWnXHQVXqyriRBTmPy6UBwNLRQzr7wfGUVnQCCfZIcw1kT/
pqIDOWGV4lqUw+R9kyEJ5Q7hNPp9718TIrDdSe1Ijk1Y0IKV6tFnUgygKKE/iYRd3k2sIqeJoHBo
4oCbYFjkSjWMSB9khJYCCalg5Ns6OK0xJvy63H0oBjLRV5LnM0Amlydf7RPI+mmbZ4LIZ929/Ity
kSSYtk/7vc6QOe9pH2Y/ifO8ZOVh+ZVo+3SW7TawTIVX4sjNZVMda2dFyvoTA4+Evet+xwmsNY+t
ioVYphLpt6OKoxYhU4cmyTgPVZGeUM6AiPulFVOTAg95rbIl/QHFfxevE15aQFAyCjr5Wwhm20KH
BbTfv5vNQbFOjlF6AttxyspxdEu/yK2GJ0dRs/TOba1QahHV68YGAndLgsNHpbErhOQVNQd0U/kh
go9rI7wgReywGk84obGanBfkiEtbIHJCxn3SukdvHkgRrHIPbMOxjMrW1Pa+Ptr7mYjZX84dMKe3
WiRc4UilAMTJNqqqBZY+racQ10Nv1WiNZKYsPQnjdNkYpHT15ji15J/hAE8TpH6k1sCaM3NQgiK2
mvPkc88dyXMK1+Pq33H4XThe8MLPTZyYwV1/1Hkg8l32QaZNOQ+4K0BOpnXLIKMVetkSRdl4Vgps
wwZGy/PbFk+yPWvLHq34Su0Vy/azYfZVweQ+WDPpNALQJzKTEyokwry/XRfU/Plo9u+cOzmG3r7r
IfNt0cxt0SVU7oljE7C8c1zLIn4EgFMpF8JHzvUPNTvD5HgO5E2UuN9jhsinsaYALT8x+wRVQjCB
kC2Yumzr477xSfT+xw+BDyJT/0aVJRiE/JKikvNO7e8wnSGrBzwMnlOmq47NrcqglMEtVo2HXCUn
66vk7mD7nqVdvV8ssmvI7WCi1vmVND30IJbZY4rTn2tunoQo7mPFm+vSkPKGvm0Sl3IVkw/m4l4x
PtSkBHtkVJQWRm+g/4KLBsX8sw1dTNOaeNpZinYNIIrWWusT24McpidVlwwSintWjuWj7v0e4rYv
+o3BtE9T1Czgf28ySLV1hyW1ctE8p1M37hhAJvvd+9QB36oSaTbXUXhyjRsr+8AQob8KOJlabIcm
IHavWaNcfeKr2VL1Lpyff9pWsqFtEdHco3aoEk5O6vz2BnHW/LiR3O8lMEsnbqvhzzglWKtcW6+Q
rRElq5DYm7s1vX0ylVG4ML9ZDJ3ZuhzCfz8/SNDXnmtz5IFpfY+Ia9bxb/FpqoQbbgmtJdYR4U4i
6WhCCvRy7df2OrQAlgCHhQzod3A3OEOlNJS4N8G8/HqnZIzXka5u5tCceks8MdNGiJtbRy0efBwc
qZHouqtJ15NJLFng9/dPCInWq/CnABdOBFW+2/6sUsfPxkqhl9JzvlemAMg0UxGhKg/rXfeeAv1Z
VdW90rdS6fqBpHJ5XA40SfTIQgct11fxVNLWcvyTwIaQ3kbqxeiu97fmTi6McJYY/4PoILyasvvf
OAckKDWRUAvAHB8Ym1kuCCsxRnqH+moDtlI+D9Lwqri7SYpK+jCQrezSLKOjDb0GeA27iDr7Mdbu
Z9cpjpT2SAh4Ig1g4tbWtPzzERF7A7TrjFpBQnl88kIeBz7eUzBk9j+6NtXtCVR7QvfU3YWClp8z
sd+cF+sk7De68Vqu2EvAKYximZy0uyvXS9L7LS/cV1LcBSy5v4Mk/4AgUmoer7sPFJirSCMcz4Vi
rMJypbNPf1rb2Spf7pkQ7M4tjmUMKaUK5w2HEbv3wgHjzaY0ZFZwozXHydR3EzgkdWVAgzRdWWdj
Nj9n6E9vUY+jiqcPqASm8G/sksh4GUtRtz0/ifO5tn4zLENRXTtmApOh363l8P34xlhiE49JQ5tY
hGxSAiq1aqJGCWfzniVt20YRN+5k7FbvPIBE4DytA2ku3zSrIx2Cg14Iq2nY/cNdnjhBSSmUs+4V
wH0ewZW10serYrUCjIlqV/R6G9Gu0orR+mZHq9FVDqxat3il7fnbRxcNbni2QOjIsRu0HlHJ4d61
am8pz2rcLRt5Flw0uS8GuHPYs3GwVPl4kTuA+ahaCQE4PJtnpArf2X7jpwzrnf7fmKLGn5qj1bJH
VESK3nNxXsgpQfkjx8WOCY7vagDgvHKQUZnrd1hn1vKlBepseHlLfLu8j/aRganhgeMcDg6LerMv
Bz3MV5O/z6r4l/zOep0d+fpF3GLJQi49jHqX3jvNGnKPXmesbNESMUEoNqcXMKsod8ntwj7sSSC6
qR/cXKYriwGQMtwV7kC9MUKwZUlI1CKm1YNdLJ8xrLv94fn2dv6l3p3a1HvhS/vvWlC27t73HgRA
lfz8OWkdgMvE7xtijhWfoJgZOLiIY5/lEoST2HUDP+wovllHikvZL1qeJNlfeu37qUcP7Bjdk/v7
W/5nxoI9KL2/kwXQeLZErjqk2ZjjeD+EogQgp8AXm3BvlOI+PhP+HhV3J7+Tl0iYsKqS+UDszcA/
4Z9MMV3H2zRHYqjCTR29CPs+59z92fPStfg1nFVj1MdHf6wQzH/OWXIyYZXZce01iTIlgDQcfE79
Ta9T9aGqRKWBxwDkaHKZWn7CD8dyl9bbf6gigDqPc2t2W1mQdI7vseisVgnn8dyfuMqcsMllIrFN
heaaTOM10SrukkPrOPINCf9T4CwikG4KigoL3OBypG2NU7uX3DMwqWErHpIEhIOFQ4T2MhGm99CV
5mV0I94AGmOR0ACaWXI5L3Ks2g7KM9SKIcBtTjCaLe89TGCLyoPsZU03DQS3N1p845XAV0uhCQ+g
Zifq9P3vVwKXCVfuGd7U+VWQXp/ocB0rcpiwtE3AtOZZka9AIriktLH75U1waEHOIcvO2FMZoBOy
eRbqWtd2zCmhEdIAqZ0YWvIaOUiOtpFEdXTXM5TFFm68IqDAu6yVrZKmbmMfexm0GawyLVeRz+qP
hoitlGFPTkOhBag2wxhTeqMGs/eyWV9SIQ9xki9g2Lt3H3noLkXzpWOszXpCelZYgEHcn3jP+kHK
wtB3ksExtQaympuuXa77fV0/r4e+DApSyxXrODwyHsF3s2vIGySGVlXzD0Lxu8sgfy6xqhSHJL+r
g89wtVTRNhuihBHBW8Ki8vytrzk4yY2RoJ0IUdL9vYr07YH5cO2pWpDYL/I8ErVZvkKXNGvKTfB2
n4rIrB595CPzP31Bbhs6eIRxgA1ogHEZUQQ06HNLlcDcePnUNyM7uUKJ1VMX0w3xrVW2UYHwJ3Cz
SOPtAEd0mLr/gePgnq9uYO5Oc9Zg5d4SNHIwm6/+XeyopINdl+8MoK5pDIEOxCMW+cg4YBPaCGJt
SKNf14pTdwdAAMscJv8Iwzcy4BE+FN+RvfXgmLT2bVxSw21EOxtwZ0aT6te8R8LcEwB0GbXmpswk
IZkmO7TuCGyJ85cD5qtR2vKk41Kx/+uzowFkqqU1rkhSXcNBccJbDequ1LBcpfXLtufe2V3+fxxG
jUSSIcTlDMC8jPUo5TuqgkXEQFneHlzVQ5IHyR20YTHyTfgi7b+GSCyfKdDx293gFwSzCkfaXMJo
xpZoPTcFxX7qmu69bXl3aSGziz+a0nGxjslt5tP8qY1IZKstHR9R8uiaT3JkZ6elDshxYpfxFJK0
sgHS19L+GV0UTdiCHrrerGWg/3Y+JzVUJvVpl0S+cyW21XinlCw4rZpzXZQTLSr/OctbhKe4eZH4
ORsn0vIRh1fBDZ2H2iXK2AvAorF/cdyIIGREv8WNOoOEqFJ1K6HejCgbuD8/KjxdKrJqy92Oe/nb
6cquJSOIJ0/H3hd/xQzB871yXBQGM6wFD21tFeAJ9cBnAtfh8XNEXQD0hbVlN0qwNdvMKcE1sIMa
NxsMW3rzkNWPSzI0DWBtB+SyJSO8eIqzKEO0wHaP6aolIjrWpCHf3WlZW/W9N4HpQpdSInX4Hvbl
m9W+lGvoN4wwHRCwtjcoE1TC52WqjqmHRuCRo25AQ6v0jZkPVnIefNQow3ROmuufldZDi+kJD2ZQ
SFWep2EdO/jVYC5wQgM1Ryd+2ZDuhILLXI9TEbXz1OZKrx3vuREy/vvbQ7x6PDPWg9KszzX1XE4v
pdWpOaxLs5ouYxdLjdj/Cstj2X9zyrBeKi/qlxqALlS/GNyF2XQnCeD3HZ/VM+Di/94AXBxFNNrn
Qc4wBBOjBobNUOsHoY+ySaCLA/FKgRO5oVliJ0wTepqkG6JlyXLYoUwLnYJG9nWNIfM+nLQa0Pxm
NL1qOfyc8rYpWBoglaxUVN5yyi6dSuuL8aFr82+ECykv0mYzeBxDs4pSltIWHk2r+DjEuisr1UK5
ND2Zw0p3G6slXeEaxvs6fmQnxfq6/CFrYRRR04jeNb0xWUL7X5Dotnnz14DOUiQ4kqJApbHEMHM+
a1BR0vd6u4CtnDDVSUy/hvFULly9PcDbjW6bgVEygbvRUsbB2SrB9OkQxwgxZxRmPLXKF+99XqEm
B32ulZ9CueTbGPhpgwiYDtwp6dtbbLwLarUaL0e8IwrTP9rvwqmqEZYN7M8f9S2Aq1z2QPz0udYg
OD3YEUw6/ujYRnbuzS2Cgu1xhV9ih2UJLuEARqtlHnJ++Q+3VGO0A1gOy/TQXvnfv2MhtGBx+L/c
JZbYGbuoo7V0TJbynRCpxLqF2PTm0CFusp4xmq9QnjNmZk2NdmGyegLjyB7A3q+ICxj8rYUW4G3/
LTCCisGnXWCyM6BxTlrU4fyJ6aapqxSinnT0KL11QrIFX3utFelQCNIAmrPMkc8b7MySB7QCoX0x
/3qhMFlhhJ5vUEq+kTRy4Z1ZQ2pXbNJb9rKtFuPe82Yku0OysAiuf8VFnjGZid/gof3/FYmW37LR
gDiBk+xbWJcko7iGVgBOf1ey1mqXsPOnG/P3qxnubwminDbxRGOD1reHQ5DWifftM1j4cSnXm8MW
IS+O9TeI/MCP3IZqYQaTSeX3x6H/Vptz32kDFsy7QPPYdnrrrXOzpfll5twdqKZMIKntjMr4ZDWR
rFz9GkixNIdmKg8iJA9CkYBxrEAbPEvvuTL5xkxIrh3EezvSlxHNyaqw2mYN25GnV6P7ozOjeU3S
GcRz8OR1ga707R0l0Rb3T0c0DqWv/cxSVREfbJpb7oZTLNbPHw95RE+3NeQWQcsCsYxE7MfzRryX
O2DueuCtTyWFqyQHk9/Y3iRBi0XMHh/HgXyP8pHhA1NfYB/B1nTydanMS89eHn9awARcTKSaXHe1
E6B6k8z0ytnWQIiGKK/st70OlY8eBCKEGbGHZhy5N3/La3HInIJv+RwGWU+2ko7jatKyGilre+lI
Q01BhjA0WpP0VDVoc32LkmoAzFii1bS4U628uVYZGnOfT0mDc7uWJcniU3J/GVFDEMv744dt+QhR
SVYUx63PcIZbpraTuGcetE4u4GgJhmhCNQPCqve1XVajL/WcU58laF4SpdpagU9fFjjVFtHSUkbu
o4bPGDwbcOiOs1aEKYZAzMKNcVWIJUxRe5f+nehSyKE3FYBZvCYnLrzg8p/W+4t5qd83zLH0vw1e
fXPjy7j+aDS4JANrr4jyMDnWQVvLfy1rUlSee2gIn/xATJrwYTiGMpU9OSwzEdLAOrRloMDMbX7p
rR2mo4XZ079TTejIJl5YEjEBb/fXD2ewJPT+C3XUrebFL0iU3R7X7xEswPCteYM62+BVBh7fUi2U
NVDwmFKDPUMG125ymXDOr0Fmf/8YHPC/PItxVoONbBmFi29+Aht/bynQwG6UGx2KDTnWpK4ZW5Vo
s1c5ezs99OuqpN966FF1A4ctp/OhkCV2iCrRxjQCw6qNx+aodwyDFFRMPRt363sclTWnIzVPRDHx
H6yStK4jl1dJ1AfwP8cSx5BEpqAqJBM/88v/WhZzEboJRpf2aJYoVePcPr3XJOJ6rSBqVDxouxtZ
ne2xtpID5OeuhrYkVu7uGJVdV+cgbpHleN0Gb1i8es4yfGQ/fhB4ZnMLIxpfYg8q9Rk7y0OZZYh7
6WYKQSe2EDeA/7zyVywWa+dTYlR4s5N0Fb5Th6n4ZJ1sXkXEXxhI4vTd/vo9kfHNWvy5MNAdlI83
lDpkqUVaTQuYvqXoO6LUGa4dEI4WXTfF5U2tZCO6OkoA8Wh2E4paYxq/oTsWJ9VZXEEYndqP7rbG
JfY2obyP0CrXWgNvAEKqiNenOOTmhiu/+jfhR5hMbLo/jpFvm5T6SHrrgy39jwY0hhGT4p0roOGc
/1qpzrqCHMp6Z56m4nuukJttXQZ9EWWWRQUXqgIMnKSPpu9hcI/rygoK957WRw0bvoZZBLV6ICGT
kAtbEr8D2WfL0exbNnOj3uFAeveDmGBvYw+XZzCG8Ml5uUHZ1bbCpcBOJbNDK76IGdMJB7WL59m9
+e2b7Qag8AJiO5pEcQ1M6G+qVfoPyISeuq2ChSYCnBOcCEH5zjernnE5SdZn8wLX0bRmkw0/iJ9p
xRdn858cBEmFezxavju3lMgJ5d/IxtedXQnqO53/AbWFAF/SgIn+4SxBybfuxjMrkRUZQQHH1y0r
uHt+O4gWAY8ZDqJdBRZm1kzc6x6YViPho1G6SMW7wvSu0a4ytsbiH4It159469k62yKe4LJAFA14
LPp3VFvRI4RMlK9+xPv8cP3/uukdnRCImQvM2Wer7/DqZHc4p/fKCoe75GqzT7C29GxLKBUj//py
7I99IDSR0KHNHTiNJtbXACX0E2Ew8MC3wciGpriEZYZVZo2b7M9v8O+lf1I0ioCeIe0FQgV1TDPW
EivzCGFLretRwncfCqnF6lxIgHcgx6aKqpa3YQTFVtUiZaos2q7LjfSOeBmmD+HsjRTGxZgN3L6J
QAk5x5HxmG2AWIhdNzGxRBRrVTDzS5e0BB9DQJ1FyAHvSAwO+rIwDe2ElFMAUy1OiLHIOVMnAvah
JX/RK1s2feLA+NqOkvgIxmbmZEMHoHdGUCdR93WtsZWRHR/bCgXyeEnet1xR+YWgrE2pUm2GuztX
jir3HQqxPX9PBwsUQsnXE0lEcTXyEqUq4bfYxc+QnlVCSDeeVioV/V5k44a1KW29dn3fNxW4SGh1
iFs3QzXoCNpOjUOwo/qad2qHBmRjMZirPcvtCmm1FpS5yU3RgCbxVyedCpVztFcJwvTFZyPjNIDK
jWDKzk+2OjD2cwhnYPRA3ynqqK5wqYdx71peXxZA/yEuZDAQGpnRGPMIXizKi13esDZLdpkfLwNi
8MS2yfkvykqYMqCh2YeW7qNZdWmhPCCnAWxJT99dJYbppGEUZMrDp3wRxug+lef5DnX4TQqvkL4y
8Ywen3oxcyMoNSgJArmVsQRJvIBnYlhw5Qx+fervhGcTfEe1f9GrMadymND2JImefdt6/DXmsQKP
mhsnnvw/qVfgMzVn38sakR9wP7JShrhgmlSJr87uECLfGbyo5FoM9VQwCZlrpXmbobKtAN//hN3k
RMcOam/uUlmz77bzNV2swYS0opLQ5UQl7IEKZRHrllV00rdm0bRNXQ7zDCkspEVNVbBUOJ4u6VJb
XfgiSvBdM5sG1DusZoMNdC3xMABB1z18z9ZQUVjmJ/WTTKMeW/MVC40DLNctvv5Ikj89fcRJHkQj
huW5HuEhHd5TY3388yc3cIJ+bMEM2IwOI64U0gV6cXCFVQ5DXBSHJmEYCJchngV9Lx/9OAhwup+W
k0Qee3aYITSTY06JlC6zN6cw84f4WP8gZR2HGa6aEBlVulIjjPDQvPuSL2SGBj4P6061wSuXblY5
lXGt1tr1kJ91gadnAl07dj47ENokvzMA+8R1ZczCl/arBWsLtPszBBtzqK1tKhTV353sMzfTfuCu
graZTM0HfjfQLq3ZuDAQvSC/KpB937VF8t2Og3cDxli+eU+xv48bZgD8X/AtdOQXheZ5d0baqyd4
ZQMydRZvqKCWuDp6Q76R2beLuOChU1DAbUI0J/fQyZEcenDx5gVhcweJNa4R9PevC6qPUdJL4BxL
1EJhfuoTea+K5MjGZkd85s7cUXoxepqMEpgkNGahb4jPUxRd5VlNUeK2b8XjCjEN3u1adw8e2ihL
FQMzI8q7lETLFA8LxcjIoyzQQqVDntLSHRi15O0IPgMz88ihgrMaKGk7gjXmfKN3GwEB1lAQfiJ9
0/w1S3utGpktgcQyM87tlY76ub2LT73zmxXFGfkMM+knuPycauoXmli/eSdvMK4VVks1Mv1QaB2I
PWJ1iai5MKdGoRBzFqzAqs1cuojiIoDWsf5iUGkmzE0itBiX2crv1hZZk9vYjXMTAkmIoHIzzjmV
c4QZOhf6Gt/KhIvZDfH0fGuIPEK+nz+k5eYNDOK+DmELrRe1yGmth87HSGMK4/EQqE3wh/OdJAoy
b9u4+ITvlFsba3rgt0tUF1oFYJ+LTjfWKy1DhvJUymsz6LKrsBgEmFWrMYWig5TEydVQHMBpY/Ex
LQpRuYVktsS7xtMxjfwWegI1HK2fClTZHd9Yz4GJqnm1Ms+8MhT1m81kil3o8oZKyWh6k82/oCZK
R1AtdB0/XWryXoDBJe1uvzq9kH73sxFmk7vIm5haLwk6OPlZDKOiPll6d2x+SfJb4xUDWchHw1Ez
F56AYCdEdIpgEDzLYpl4IRcsUzu4jj5URNXETUk/VI1B2pFWcIbxmdFco34GDIu3yyVDYqWxOA4m
Rad6bFm12vTuW8tzhicfCRk0R16TFj5bGfwS/c+xnPv5I6HKg+v511TpNrdOHT/jt9M8nfSIP6u1
RiQ9yp0Fn+EemmR/n4jYYgDDJ/0ttGv7ZL5YQJ1Bgt2xX9a6oRr5oW/0miuO3nUz12+hJQER2J3Y
2/wxK0qvswh1PzZ8OJY6K/L5VjZgQA9yIwkMzhA8ThIkIRNG/IKAvuJwnDdel1Yl7XHDUtMvENwG
6iISC2+3SKbQ5u+8Zq49kk1GPfvSQa9iz8lbzaTu1WouylSGCBj3xFwPf6MixY+PbDwqcmNZe7p6
cXuex26w0yBtJJRQDY78YckEHGD6f395fQ28N0V2zuN8CWYGEIiiENkhMkj6ls2HkUOXlziQTOJG
gN5NEj3dCqC9l4CK3Te9gS1Rt4Th/sBQh84UAhEJt6GO7fBSFkHe0+vKdRdRDhVbgHddoxD+rpCU
eSHxM62WrYzGbcDYpfm1Xabtl9QE2t1nv/x2auSpBnJ0WgPsyoBQDZa9PCXc3v3iJ2nwnMOlBLln
+nKIQ/D8U54uyBw4LfpV847cI3MSA7gfEyflgSWw3FGircryFhIV+YVamf0d2HoMoH5Skyz8peuy
TZvmy0V0mjLU64GRIJMsnaUfyCqXeQcscpBfDPz5cp2mVcJLLXjblVimFzkVUcV+SXfd2mGfcbx/
hSLYuz/8c6hhF5eT/4/Q5/g5cLxrLptNILCaybnXeFHu1PX/WorhQ82dSakRCklU7KniNq50TCyI
4SF6DLoXC5q7yGWs9WmWG8TVSLEio7Yfs38KUKilWqHuFrwI6NGeLMbRoEo4ePLzU638oAy/FgYC
w/NPYlZGzOeoECABf7xiQ8TE4xaIPSCwVLsQUT6NRoN6e7fPCVT9okaaWNq0omfX2BIPMcX911/i
HMiHVD9eCNNTZAETtdSJ2oXuUWxVw8ZYw0qD89QN6AiBMuQ43tKczZgTgdboclHmY4LFYrdGJcLv
k2WCVl3kzVRW8UcCVs4jnOrlF8jgh11j9FS6aeb+XJVj9cvQD8l3TSaxXJTwClQJFRcmDBKu4cUR
OXJ/EsjuHa43Inrx03LOC4C726jkFegBnwFk3rysIn9jNo6rB231ZpI7Bhnji4+c8CRXp8/lVp43
3y2C2Kz0GlYGXYKkL0kSKibrQHELHmkGYiVXtytNhLwWpQL6HhNNJuJi4FcnfeG2tzr6OJ4oCkLy
GnfY2oFbd77YA2REZspm95TK3K8aK82RipmXBQMPf76EyYVaXodnnVyRydo3lnQp589u5OYUb19V
HjDgKbLjIOJFnU5DYHA82Z78KWnCYw3d0aU7Z5CZQlr1/xTxzQ16JueE3jokYRISXcsOh2XIaP9T
RBpm+13z9TM2cDVlOLXcVaN4Dj2QLrKh1mRxFLMKjklvsFA8OCR406QyH9ov2ycSSwCYurQ4l7cD
3ys3Lu7qUa30abQBKJXtvZJCP8F8tk7QUig8lMytpn0Ub9vT6JsD1xAx3IFgeCfkp3N+SlO0MswL
/m4PXsGZo0oDxM5UFP4ybbCMaVqrtmyy+Blekxg68wNRjo+MMuLffyOkmNZ5frcDHjxsxqgYWP4C
JoWzBoskcVNjQGDGTcOYpBqsodC3jQIK3qQ6RBaNnT6z+x9OPcQF2C+p7hINwpCEoo/sa5jAvYNq
mSwAxPjf44+rE45DuqPIluriFRP3bHvdB+c33fbOxtoWhHFUGRRA4WawBGihIaSiNQFruUMQKnqu
5CryolEybkPPB/GsirB7e8c0pPKwU64UNz1SBoV0rtz8oXHUkj/frezLZz7BqfassWSxGZJr0NSm
QLA8eihh1EeGMl447DzXaFl16XtP/SAM4VUXJoscUogATUPtZR3HElLC5OxQOozrxTl+wpdxfot5
iIfK+3fZ1jUjyEjDG+Ea1ZIgqoV5r0d5NuMjRMdI4FJ0FKWHdQmpd7ziutwHCTudpV/b1MQOs/bO
+g2jwUJgeV9Ij5zSybHGXMvQPdGX3liJrPzp2IgIbQGHN1jm4xyD+9rr5zJHQfXVvmHTCAEGj5oy
lpUMlXRMFzXUZ6vTmL+D9A30Wac908DGPseA2SCBu2ZVjYwPixq+YDBeP/3nMpj+IGkkhvwQMkTj
/o5Pvl1tuN5xZbCkPhWtmRDhRyx5tLBh9JS5hB9RP46Wj1/EzwUP1hvCS2h2iC5xRmJGOEI6GnVA
Y7akGWRHC7RDl4eHkb+waQSRaiyIX2gytIsm9WHT/0NWZssMr6+Gdq6yIle/pav9wRH1xSiMDtDt
ijOu+soJp209wVWhM0Tr6pMewYU796xcr20CV138lwLp9w31hcNBxyGgzkGRxazW7qIhJhoA4woA
SIKdT7/neVdSJ6j9vokeKq4JMYtgr9g0s829AnSLW2M2GQ0GliuUuPCoLSCBa0vjSx+LqFFa6hR/
+GnWmJd4Lde/3bOn71Sh6cdM5rUTfiD40yVep4n3Ta+KXJo1P3cxTBoUeRef+9h1tTqDtxKwHZTN
nq9Ke/YwLBO8akgXWvr96EBINCCu6RCTV67kmOynmRyIq5TNMhFOtoUo2xuaZb/HBklYbGBYly6c
oCMgAMKkJ/DWrtNaJbY4MUhjuzMp4qECSUJFHj56VSq+n4c4FEY5HzJSTjpBDpg+Y4jHTJes9sc9
CtEMZwQG5SAj7mooh50fVAfEdAJJ0spywxCTiXIDFnrFlTQDe/kDc8DsNCPMKJCVL7DwPWudK4RW
I1D4e9YwaZ5XJU5NY8oRfSswhTxbyaIyFd1XBEMpmJfZiS2hV6LYEgxEsLpJuFbj+LZFpsp/BJx9
a4Z4h1mMV1g+ek55zWKQoed+krVkoImrPLOoygqob/MorlfFLqsWlaxd7V31AzBKTbcEbvNcu+iS
1zQTz7ZOLf7t45UtRwRAMEk7IKYNWFqWtyAjnr3imwqx0Hu7ZeFK3awTnceiQjGYVMkKQBtF0M/d
HAWdIluvXsc2PuT6/H1lVUrgRcOMOzaQm+Uny2MdSUGtZB0J6txXE3JyJ4IuCE6gy6NiNOulrzoY
kKhsy3Bzs4qV/OE5WRYmS0hin6jJGHtpIHYSuWhLrx47iqR7oizKF2PXdm9F3TiDDPNh//e06Nkt
R9MsqKs7UYvaL7Ba8HByzrcIv2e9WGRrxqb5NneMhgUv1rVD6vdm7l1iGMOCumLA4AEY2lL5h4F5
LMGgS/0z1eUg3AcGJ4jOWRYPi9S3XlJ51f3S0ZLCn24nf1UYZWnfdKO/wW/mWFyzlB01u6Yv19ym
mDboY2oKxvgCWw58Zf2JW33G9+kRpbzPkDMaljrHDjgH0C/fWdrA+GbjU078qfMhDBlJGamq2Ltu
EWndg+62RRX1Ga7cY9q1Fwi2oJe1joWgMAlVJ+o6cuy2rRCPlER+Pvy0c/VdOG90CXti8tH503a0
wXS2B18HyGMyx6/wgSUC2OUVlcGBfSmKJ9Q6BRSWlh4LSKaHYJnnDEKaX06v4QXQGEEXlt152eiu
X6waYDiVLqV4Er4Adawjw26fw9onMYS0ECaFpGB3/Ek5pJ4eTmv1HwKJSV2Spp9pfzYi35RlH+fD
Shd58U5HX+K2K2tOXTyH+kiaWGdrCyC28D+Th/WwfihwgXMQQ93yyXjcui0J4d0lEfxK+NB2MU7B
uNsdiMe10J7Y+lnHFlHD9Nq5O/SBt0sCNiBMrqVmfqEbiJZKWiXVy56EcGsmuHAc5/es0dGmE613
GPPNH7aV3AkiM49N8DBrOCtsNFt4khWf4C3TevEXSkXagLGDYlGyvTSxPbwRTZufpJ8dzW4lHWw8
SJW17T+xZyzNHD45pZUd0MhCR4BuZma04ExpI7cpPS5s/u/J3Zvigh/qXA0GoT/kieSQFLTnQeBC
eAItihNbRbCTKnHCl8lGSTLj9ls+HfkMjPZ5+AJQzSdF/2lsbMQR5wz/bvDdsjPqiPWeRj0P1xe+
zfLZyqCDp4N4fR/rPOA/hQqe7ggcOe8T/dzLb7yZm9XadL+xMfughMfB7e/wL24uHoDaLv3ujkVj
zbgud53scBT1evPwGKgL0VzEwMfU7cjJ+kXfoF/9fviIyV8cq7oRTpchIsyE2axY0A0NregEf8b5
6dsqi/ShXhtf8eH2/TmOftJrjapKjDPRvGwr7Cgq5IGBDgKE5LFcSA5A3g2sG4rC1Nlf3RhGjNDT
nHG8VQQWbpGRnaM0+r9abV9bIsDcnH6QZm6x6NtsJVZNIsNTzNP22R40/CRGKPOyem7BK90yEmqw
dkw1xTYpQbM2i4ygDLJOIgF75d8s+21Ss1s6eTvI8r89OCgoVWyWO4PBVKWr9y+Vx4uuSQl7mQui
iS3ywuRuxwMBWRk45FSdZp3Zjq/SlXyBZXO5Nv+CziILkTRtu3+oAkfif+O/YCImnCatHyNtXSgh
CgMNA8UzF7dpAquO6LHBnR2QhtU73RmByoxzQKPUyzJe8MwduDFQaeNZVcPnwqbMs9S6JFt2saLx
Z8Ms1Vh6rv3Jz6jkAnfYklnRNGcYadZj0VAkOOoU4VpgrsaVJEoeDqnkDf9aJ18FlLH5/GvNdLFv
SuFycQkFm9us6wISc+iRpY+uZqlkkqz60v+G8iz8R0wEJB+YhKwikpVtqXP4rxp1nEEWb1DtNoBV
keByoCsx21WWINnucZfVWTmL3BozfnAAvymm678lrnQeQFwzWJMEN2RNzUwmpuAAb5muO/XyUKiu
uaR0JSTXjRCmRhELs953Gclo9n9IHdzrhX9ScFb59tp6v5Ia22QeIpRbqOy636QzqXBiuWucJMgz
vk222GIWlydySyURi2ni4lJYVjOUhkdth5HV+tNgCe9h5gMclUn/NxSp6c+bemyWSqDtqsZA4dWS
xrkG4BkAhJdDD8SGMrsFrnewuTNLLZk8vGq5X/0u9Pr1cNdLYYheU5U0av+QPNsNw/XLt6AE/U3V
epk9bCcrSLOHHHDfMC2SlzdFp70VXlCd3zH6mQrXfH3ZsFQReXCDuqZ83zIacLTpRDRYAwAbRCFb
jF1Pg4b2fJkGeEgaiFGCszI3WfLS/p9JTI1xdAi1xnTc+MbK3LG2bf0kT99nafd/RF/8ssk5a3e2
zH5eHl3Sk+oZ8EOxvVDNFZizKbwGt9zTtTMpv8ZPoTvYUETdQfHcMEcLt+0TF+iHqpZO8oWXs8/L
xI9+Pe01uNCAkGIX1F0ghyJ1B0G55vHKkwgGLWjGMwOB1fKO2nYlAK2oVejwKAzpnfhMjYtwNs2q
ViSmLMClrX1BQhUd/zihwMhW57pfSMckAOeJ5I7yR1e+00G9EZpa4RCit4lmWthEZ4gL0fBrL21S
ieew2M1W4HXwz5jbv55GsDLEaaoTvgLZ5+prT7ixHS4cbHL0A9RNC5Zl8IpsaAjGJTvgHrmj3fST
YH2XXPPkUnaAImit5CGDUCpTeYVjccalB0tkV9dBlLhpuSmqSjxF8EZs55pp2zotTOmg5CPwACNx
D8J/Z9mUuaSa3Xt3RLsOrI5qsHX6OSM0qlS2jaupXxPXOz3oV39vx63Vz1G1dHSj/GcK9hapvaS+
9Fai8CgkoX6yAK88OxzwOZRwq71G5jKZYh0ytIPhfQ7l+1WuqFw30uGC832Mr8hPhJtXE6Yjw/1N
PWB47j+4UNjQSiVfviNZJnMDhPDzva/3cqdgdzChFhQTyp3kpFcdLGm9bbz2modvBKge7Hxe//WW
JVBC9vgU2OsjfIebbXFBd3R/W+1e8asUNSfx5DtxM7tRObOaKhX6nbMV9sxZUzl9Df8sUjhGHb4j
zBuIeE6ob4mRoL8ujlYB622jrCZNS4G8iSewKnzTgmmlpuo0dh45auz+dyKMPX8J6pC3l5ccLNlx
dkILPENcihCa2r27bnjEMMvWoYLLklKXbfsz4XHVXOVZjSbjJdleDbN1D5So7bKB7mLON99qcF5m
FE2U0hNRvE6JZb3OVAgz8ERvtu3zeUlWJDHjaWLdHTL3gubyRoDNPNTMwHovTNlGToCsZoL70Grg
rXHWKSO+8Z65nSH+uG2qqV2Qa9hDZarduIReRHLjzPaELgwpCLxjXeqS3NhCiz8FIqxeayMet00f
cvGLQhxaZvaY+iZAPx6tnzKr51GIhLcVdHy7ZvIH5dibNh+4B32WgYyfBF6rbcO71zz4Pyav32Lj
2ADBBJsoJIk2bNKc3OlmK+yLz83dXtNK1OmQLa4Jux05b/diBEC1eaeYSxdwn7WhRyeJXmvKXPmr
oelTNAgDmfeuNCtYYyrt8zQuOszlCFbr3AlAn0trHB2XVahuJMFmZkg7dqCvsMiBLyLmBrZoWR+y
ZND2iA30+McW5/2UCgyFZoi4ifR4//Jo2JYZphxLhcTbMI2gOBjyWZNQ5uwJVgIuEFX9+3a3ZsJs
rkVs8WeR0Y1XBjUN2wnU0gozpNpPgBVZxdCYfD0sUblRzGyzeo6O/sjKzT3hAwiXDKJRVcd2MkoC
Wv6HRrROVQmd7uIcPamMvmnWf8+ekcfi2SyYnZ6MpnlpxWLSW79Udzxn1ipJA4vHqQfkRfY0UT+G
uz9cGIS8tyaesSn6BW3CLnl2pnzbRkqHcDO6RkquA67bxcU/45U/u8A4vHAr70kHQKEgulOmkxRH
vbETYwFKbn14vMSj+b5MawNjlcBS+aobQaTlWowZQLPovOCLMo/4uowort5SHfjYknJUpn71R3Yy
kmbsAFRxL3ktsuIC5dC9GLkEXMwqaRqDMFhTGF+6mKMhWvbthnUt7faycXbcJJBEwLTrNziNMd/u
rEgcrKw2LyVc4eQECyrWgwc5h3/cO2vVs5Ab3/FzR2WWo4aSPm9g8YmkiMZYF4qCRRNUULhlirGX
KKG2jL3Sa/5be/Vh5fQjAcKpu4B3V4+LpK2658ZMdPUy1buYoPVyVt6RZZzt6rpEB7dDd0ejPZ15
7VsRr15kzwfSeGSB0xSSZtovZn1BX7NFw3AEisrejzLSJJ2eYuRN6PWiN4w9P49yoD2A/fH8tQK2
S6TOChpUYL4OCOSHZXaqeV+HuqKTHzpZDnM6MwiFLbvlopip1ArcCvoM0px4iLfggORn/L80sYgc
UINwf8Pw8r4ta6Ny+3P1G+xYKsTTScjHdLJUVOqyKHl/z5VP/ZaDRyKWl2jf97TOHl7cMODlEZhF
tWhXMGmjy2fFFdM88y4HU/+HdqCu35PrHtXu2yhFECVaNcta/Vq15slh9latMCN20/Rc33Wcy6Ml
qJ50PtMvQ2ZQ2HUsnONGBdIrEu1f4NCEf3beeZ666FHRlWbYa0dBrtGX4UuQPD28cxtwJHEmJ58i
YN0hnMBhHZu2Hsw3AZtZjdWhGqJPY/3rote5Xh1+29pwutbWgsIa+70nv87OvKYi6L9lhvN02g7f
SV5CmCdSY4HK9Y2x+YVqhSJ7CW8E/QKR7KOtNYum8OJTv5QAWPcjEomPnD3IFHFGDHKZFCZ5bfgu
mGOtV+/OuyOrfWEReNdC5hAHmGVobG0feDw668/LAjNW7Zyoj3ctv13CAqO6Pr9JRb8/aoaJOXRI
Cwi1rk0j/YJFjeexmE0s4PDLQhNXqokk1dK2/YObt+IrfmowJ7N3j1XpAGQ8f/x7q/E9YdQDJUuy
21MLk9K4R/oG768//Tg4n3b4OpGjrXA92f+uFAGnQr2H3nM5f+J40pJ1ixmZWyepUnD+N2sYcKt/
fGbZxHK/muhw/FYVquK7O5J8oPbGrX+2BCi/tETz95lggj+OcDdr7z3XG/vtQPB4L4Hp0uV3HmEy
KkyIKprsrcPfdeJF1U5fWiLYQ4+vCHUvOlb8XjYaV4DE1jYqubG++GDCM6ZmqOnwJB+72QOj3nKu
a6hYgRMCBmULbmrO4oKt0KbZqQwHO82VAJQM6eSSlcPv+xDPVpGf6eQmJ7KvoKvUpLr/0bjU0GFF
nNnK0uXeh5d+tNW38DmPEOXix29N53qUka67slpes63UwoCtUXG+kG7eDOxs9VZPKMk/KgNGFqm2
ST1wCLOKJRMxHOF+WmqGSyZmqw7IMwMuUeCG9u8vt5s1Uqqs6n5VjHXds1HYSZNZ05LBn8KVDy3n
zRm29axE88DFZfUXtkK8M2wKum7MccI2r3E83S3cti1ou/z0ONcAsCNKsazjEE/TYErggorzPn1f
r/annbgkBVd5u1cma2Z8bNrkgzEc4Pyure08Cu+wx76dPBN9tHlQPQLZlYeTWajxLPT7oeA7Fizw
XetIui7hwcq6GNNVn/6XZIAMpdcXwrD1WqkaCfymQpbfBV90kp8oDcsfa5O0+CCEyApGJsXqEHEb
q4q0fu7khxE/5ZwbudgSe0W+nGS+TZvhr5ucUlEps140gkN3ehQwIgHL9MYLYtlU71Jjzo4L6F0U
fmVnHMfBaft4CNuW+3IR2N/qodZR6hXXaxQdCXe339T621t7b97Ejr0GRLN56edddE3lBLAj33s1
Jd71utoRMrvNdSgOUlOAo930MvJYPfcP7ILwQmC3XFtW7tBv21pxHQ1+dObvQcL2vhi4LY16hMSt
owDtwPJvi2+EHq61hyXthVfGaPYmxxnLVni5/O9KOKddB8sSU0YU7XOlbgtfxjrwgE/h9Z0RdVs0
gHv0LPNB8QDenKSYmQwq3l/iojEt50OaLPG82yuXO74iWnlcn7uvfct2mLpvXR+VO23tU4GVxGf3
fogKbDJnh2SFu6LnVmnVuhHjft7QPJicNTY3bKkGml4nzQGZROKW01Il1mteyLWGd1hv1At75HAm
iTK4R4DXC+SYDJyYCIKP8VChYdBMEAYPybD9znI2d2YHrEGQS6Fyv1YOit4+fv0Znt/sWNAOQ/74
Y2aP0MfGXUUXfEwTthmy/t16YlLBhl1vI2QoHOiiXvGiqVmGJQxJ1PeQRzyrqr/k0FlBe1TB+DT6
HbA8u2tM4TFqNLQbf0bORIfp7rsVNTT99Kv61ovy9XKxSOcbX+FNefZwIa7uUo0z8je26RCUVrX/
78g4oPkrEhHjiQcBANeebnn9gg7LgPyH1NrB2SosWICKiNtCPnQcJQnKEP7/MFOmsOuVk7TM1Z9b
RRupCtHbVGa3Rofhqd0vd9wV3KFiNHfTRvO9DJoo/K1mNKqnc+dNp9bPrKRXRUpOIqaY6kNWq+Xe
m0d86gc1YpHEKt+H0EsSNljLXq13dBIvNlPEY3zP2vCdSmS6ckjT8amw9WGnm2YQFAU+aeWM+Qt2
wbNc6CpOS7lMrzMIhXrvOEBeVvOduulQ24BW4biJf/4WLX6hoktHfLARMJcsVvzxoSTxE5QnxIjT
sPF10x6S+lCPaSeWvKgqIf45lPc5IQ/aNjFivYQpSL9nGK7KxJmYvkmO3h+mdUokuESk5Jr05ves
pHNk4c7pIJPvUJnHK+gylndYNj5Lb1rTH7vNqputc5spVlraDgGM4/dUS6q9/NncCFEo2lBvJPvt
go31xsKgFPBAEoCWEMuP0zPlLv32lzHxnJEAArtkmkPPerBNKw04C0OTbOodLIgYlZ+4f/4En/1B
83MR6O+OSTOokfvFOihPY+fvhN/MBDFJ2bRHucSJqb5zXAIbDI2l7M3D47C9TCsmHTHFodUK++7J
q92bmMoJ2amUh/t+tA+4LEFOdgZlgLTAGucXk0egspg4w7een0HkWzvLaZNkjjDPGbBVJjFxIyYg
Sz/pUj6jqzGBc2Txkpebwd1F6P5P2uCh9q0UEgN2se5jXW/X7Bb31Ap2o8nIk5M+rBu6ydnatHb4
D/h8tMXAQpKqPVJHhJBGgPUI7BVWTdLTl4/JJzugZrLw1TfPNNe9pxy9nlt2Dmx0BdZqhLGrNOOq
bYwCPCDJI8r+4bHfUeGRvHQSrMq72IeDVwhT9E+jW5ihBfqQx7N//ZT5fIt80DOY0TKdduClPgxN
VMEKnql7a4x1ZkWldyqfr+t6YuheWI+PM+UqdtvgMWWydsH2j8pFh5Q43wpDD2IbLrPhdvB9FHui
hBYtPRKmp0h2xcbaE9GuT2h/YBImMzrwGlN3o/U5y9vwXdvLxxiW/EacVT3eyvp8KfBAsf842IgJ
p1n/vet26HBVEsUlEuemkO1cnwBP4DxWGK8dHy6TMReVSKzoaNl1HoJQVEhTqcUFkif1YzP29M3O
GW1yLPXPo3d2xcIApREtNkxDtF6viEkxH8VYEJGtKCd0LAvg2/eClPnI5d5UnoVXB7ZWVWjw5Z7N
jE9nZ3EJeCtJPf/XHWVv9LEGRrmqnqjUxi0Y17sx3RYpIdPMsPh9kkTvH8+7LIqGoO6c+VtZ4CSM
x2CJWMzBvrc0z3IE6dMGcyEpNlC9oRDNLN3ARIRnV9NEc2BDAYzOduArP4V2Tx3YFoFaQ3FI3c0H
IG2lyIfOCLHaSMSKYh8R1iJTgPmqq7S1HmV2JFvilpBZVwSJmO79Tcm05wTrjJ5Ui868SbWZam2Q
L+YMXwgoH4p8YzhZgewnpkXZjaCzeDTyPUq3K6CVdr92wKDylzBpvBSrBN+CjeuP0VbxxbHztJg4
RjVha+E34jm6LRE+a16YZ5/mvBRl3MUh7nkzRlI4/ZpD8qTaa7A3l/hKigLJ28Vv9dPeepTOLx2b
IpKzjZ2FLScGOHX5TGNHQa7+Ie3di2gMe54ZpzhsYRFEWxWArfJMGMOsZ01dSY23bSzupwXws8+l
jCJCP2sMcpYCsREC0J3eDh5cDh2CbAMLNzpTl4spwbU9zZy7cO9Vdn+o5zyFMCbds42uHgwy5XQt
NxbFPQJ26UPbGxPnA8b4n4L+kTlUZhzRzdOz2EKdxZ7lhWMhztg5Aej1diZbBSKG+tZvjL6z6OLw
BZ09Kd3ao8WjI0TJulwD4SiRx6J7wMuL/1LcPT3UJ9c9qsy4vZjLgUeaebJfmBQ2wkcU3jEYm1rM
1uJCZcGyKzZOp6Ee36Pm7DY22nksB/lfLqV3ill7n37h8ouZppSpATbMIYx7GgCOREDqAqrCbcYZ
GQIf7TngwrEReYP7DL9xLmHqKgzFEvcqM1XsR890wLvvQrdR6hATTtpmvNUPZ39kyPUKvnpF8Fnc
5dGdIG7y1SzNMK0PbtcXVxktl5nzCnc4sLn6cODYGIx21YWce/Xh1ZNfftaROvgHMWJaxXtlaDM8
3o8+ocHTrDOfmD/WQosh04Dt6agE7WDY6MN9W623AL/Oz9qXqV0Z8reyAHTBhux8Askt5lc3U6+5
SuPg0EFmigx8PClp/DSJnq59OlEchgQy7uudIVbmepisCd9uiXmKYgjd/bS5b2J9lgyeQoqFxGXw
UZmkb8rmjfWx1Z3h7tALZzd6EwOOsipYxobqx9vDRDQIA4b0mp7GHW3E6CK6lY4MhB7w3ww4xe+o
tPpjAHAl84MPIUbyhQobvtnHH0bTaKkIY2jo8uLSydUAeSR31ZX2V7QsdNGU2Crnnv+xrsm9Enob
nh5VhZNA7dB35OX06HpCszURvZCYsGGaFKAyIDVd0WLkYhp0pzu4f+wrUhcj9VPDUBCutrQNN6jP
NBqNTCFzG2A4KapEjj140SGOilNWShBc37HnEzDmf/ywN5AucwKZ4sWqau4S703KG2dYk92fT3i0
aSSIArWzOe4xVyElaU+HYHi78kloD9/YRhfrs9rgrDpcbXERxkCvwGDyc1KFJO8O+rm/SPxsq/23
z21Bxpxxc9Bg5gTEJ0WFKjGUVlvEHhnzZHmM09mV6SlPSZ2GH8MsHBbqUs0J7w0cMFaC1DZH8V/X
LnKjebj62yUocRXc3qRSnkCTkoAgZL+lRGCKUaSgQ2XE8QoIq+3ApaxAq48U3S7Qdm1MeOXTy6bB
J2w4c+qhitWjHD3v08rat4LmLi2bMunFY6JuZMfytD2ZuZX/l8rTFxrsiIPkUJEmok7YeIJ5Qg5G
QJiFeMklFz0/UwNfFVYhn3TRsL+esviKUtx/7kQcf54v0avvThiaVi+DR5c8oC+LfMF+QyxyZ7dU
3qGULm+ZLAbVo1dpo3aBZYxAM+jtxwvxkhHs5e6Sd4o49Z0TgjvmbG6srznad0jFU8Ecv1i5WAZQ
xP5qHYjT/1jpv2CgmbmILZk1Ey1ERUOPQdJzO8U44H/gwUEkdLFE/K6I6pwCqW3wTD6cTw7j5tk/
bzFSpNwaWmLAKvMAcTb0Y0E5DvO9A30WtyzByZypU37zBI0hfKkqOioAjQugrbeWI3tB1wH9f/qi
swzl+whtwFLo5npgfBhhRzqP5zxoLQnTc0osLpDV4Pxdu7W+UblBbR63QMQO5BP+skYghaFfTev8
P4a1M29xyjhOVpuDHcVpZcE9FW+3fzEHRDx6+/AMsAj49iVkGdCyrvLGDumXYNBT+fvqnxMJMs0m
RRjsoVL7r+NJo2rSfRRlJo9fn/V3fhoWo2piXfmsfu/mGidnPPFkBSHsT08bP3qfsu/4asJEbyVI
3K8VIP1JgLGQ+Y4sUOFohq3//6RAzhma4EU8CVC6VYVb3Ozn0Ihyt/kPT7MiTBsLm1Dr32UfWols
RLqIChszCxbrRx522RDJC84+ze3HdyOPCq3qmjTO+hiXggK+A0YElczHluRwNFFANwvu+Q2Iz1W1
paU1G8oaVbi6Plk/1cM9jGpLcUo9x8VAMt5VLx5OvQDYQ87VBs4tkxm8Aw8AOyasg4YtaloEaiAE
/clddzNlS9sQsQIqAKZ5IVvQ/+m5ZFosGPXk9t4AD7xxLuY3v6CHRV2IvAZqpRTdeMoEty5L1YKZ
1J5HJ9Ld0SYPXYF/G0oFoRgu5KSCsxfCcvpdUG2JqQ1Y9+zXPEMzEFoddGAFLLU/P3KfPffCCUdL
EqwZvWuwrXyqyFp747vnNduIfyFQBDvMJrTpkPV3zE9EeFJEx1psTaymWHjppwc13wGnv7Fp1YnZ
HvOep4McJMXiA+taCDiBvk0uWF1qRezS/ooSeDXayOj1n17FeDwzwk3+neZQYkmOH2dhrnRwXMLH
blq9sHoJR7YJJRE7UuMpwwUy0/hvmZXVTpKlK9E9DXcp++r4xEkkvxHVXjAk1/r3a0N/zvzF/+K1
VwMuIgzDMujm4ggyLTsgKuiR6s68sv49gUq2ZCizSayXm9qOBMtEx1wk7Np6BDqs8NGkmsZrOvSN
FFKJwWIvCn0SHjukfINXiu3j93Mfr9sEmjbMpy194AH3aOvOHMdTO7UAKi5dgC+DZUUkzdQyGGn2
jBl7wsZe0nD2B4DzGW9Tkln9q7FvE5NfPkOr6ta2K88vPGksXVor9X4CTxmrK704zHZSUhC21zWL
ezaup6vQYurZCPcOiN6NvSie0axU5TPG2bqVODDFbD6snOXCYw8DFYPI97yM+Jqc4FTppmoekx6a
dnt6EEDp3JjpY7AR1YkZscHfVcm/jemKduA/zSzwyREVtkNU6BSr5kvUNa6Aco3iqdtPM9R1UD+u
cOw5F+IrVs/DAgqR2RN5T5oJfVegNLSIxDT8/39u2WrIDnIOzCNP9yvV6Gb+prZiNaHvTiXS3u2i
xmDshzs3sbIBMDkaye4A79wQaDGXp5/wXlD0dPm1xZPeF+vS7QYGWbV4NRECBLz2g70u1e1QTecd
bMnwm5TnV78YtHdqx9qXqz/LF2rUB8MPDP2p8spqNav26gcG5w+D1qgnF7yvEaFS99w/9GYJ7smn
mqGWb5U8cj7UrN9sFd0aNqBtOoG4b7C+tjaSbibAfm+U2ggASJpBhH8LHIFdLDYGVNNOH6wd1DZR
nhKhyOtb/UjHFhpDNbhmeT7IjO6dr0cAov5UHZjAKT3VSGjxERVDMNe3ZbNF0FB8ZNogs2o2pZsT
3cPNedkwsTXqU3nMegTjI2DWGFSjHuZCzQPrJ4+Qcpv06BCPETlwk9YqQ5/ycX/Ecehp86nOZtTR
0IFSKj61CInjtPtmqFMaGN/ewivrFIpatr3CHwUMU3iA+1nMZOxB+pNFeyzMBUmCjItaCd4TkQt8
mARX6whajOkpakCXv8Wauz4t8K0IS5oV21OftOlPlPowRoqp4bqHKuA40co8jV0fsklBd13d/lpI
NvDUkU2Cuen7y9MXfVtzu/oVMTEQwo4ZMpWWngE4Ynxi+HMwJixxXJb1x7x4q9LXBkkJUVIHEIMY
lywnvhJPQA9pAzuUrY4SL3x11RVwceknDdTwUZ4skN2oef4nDGXrxnEzQBI9m9Kq9YYqC+jC0XYx
s6CttX8S4SE1T/FZlqYOEd0VR/qPtrHUg9UQlw8GhiAxbuaZ71fnyPc+nLrKkEjvptGh0k3JrBYo
WcoYykOgHW8wv0Fb7ofVZc1TEOe76qmYUuZhhkr2GIB0F/yPu1sp3CxoaVhBNPAbt1/ooRmBcwjC
jYMdWlldrNohyRZejr6x1A5m858ZlchLsVdxT5cjjtL73JfR0AJ40Z7iP5n3I6QZ4I5E59PHec9J
bbt1tizodOMeVaEXWykJhTCPL70U+oyFZli+SwAJsjPZAKhWup/M91Am4EocWL3GQBxwyq0x6r6r
vtQysVZ32tJnnXiB7WoID59JOICdOqwrZvluA5YgUBauoZJV6vPiqCDF6AKDbiHyMWR6lN1WoxVZ
oeu82m+250C89XjCJRX1MTwOatKizLm1bGZE5Bzmg14YW6w5Rg+Os8yVxzQvj/GlIkfRL8YFow6P
R0Zi1PFYycRhtf87PmmCORP22ehbOFQ6aF3ozXBqKC0c6cMzezyma4IJXtCLDGYyErGTdiS6HSL1
su1g+zc3sZ68yD82K7sCC2gUNZK8Z00/lDhnGpDHZxvF+5GtZVcH8Sk5umb3lGvAq4YhP2IPRtaI
Gd7ltmpj6xSL6JNJlaSLqNX9zqmziSqya+ZerNuRK1mjxF05GHWN/YBVZXMyf4arf0UCLEsqaJSF
6nIa7w4h/NkPKe/q8HCT9v/rBbBKMdfrb7qQnZvvhCM0TUiiAmXDBChQLm1Vdded0nJkHK6ZcLIZ
k/ckODmdvqr37x2cdcLu2yprP7lOcexinAh4pQYXalVQFwpWkFJCVqkitY8wLhjW5UmXMXBKJgWU
f/mqlFnGQDul2YownAOyqqF0Q5qCVsNRNgHR4JYfaHw9EnMas2QJimank1HRsdncKdt/Zwv4oHwQ
tihFMKxnZXIWZB2K6G7wtEBba1fhR8p5o1JiVcdcld8hUmsA52xYL2tN9zSGph3XCJzUlV+2qOIn
Qfc7brK7PYWMldQSbLS6WcVZc5GQtmF0g/n07XNgxSaFf9e229Ja8XlVeFSgQjQFCJcTgzP5fIsi
dAPC8TQfBkECI8aKe5z8iBSDKWHag+gFLhRiU2DElKOcH3Y/I+xkEccXW+x6yGx8rA==
`pragma protect end_protected

