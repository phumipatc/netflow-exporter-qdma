`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SWKIgeMJG6ImnhojZml3UWUckeHSRJ8DVIgQGHfd8qgDJt3/mSoKWtHTNhsJkhan15B1dShei0hG
emnn7T7CH+9sWE8VEcjhXdqIIm095OiePEExe9spXU1DLHgLE86mdF7VVJ2Q6L4UE/sYZZpDV4wq
TvupKjyoxOEjxEW7u350EUktXtATO3PfMYGMcL/2nflMK6K++80zlkE6znz/h1ptEPjzEzxK7P6M
fBvVfPKgN+G5jMkOk0llSTLSOqzokc3fDxQd2VxlNOKPIkO29fe3ZCCUMOfgvQudoJx0WX6O7ICC
oiDr0pTvenioEamakbm1AoN4XwL+vJ0wxCW5dA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
Zc3R88+67MPuaRV3MHMNfA3BaTncWPfX+PIN/t6gJoCNQVZqjA6KtTxOaYJnvEfNzoPlc+7yUzMN
OanNKF5crBDn2EEUOicMWudHI4+HzqtfSR9z6RfLZEGaka/oDGK426YqebB0qOf+DmUoGFmy3Q5Z
SU+shg/e4ibqOjHLr/maFuTPK+0VHU6l/uzq+XEsvyC9CeA4MsvMlyjrmmNSH2bhAL/pOQOa4749
xw8w6Uv76Gpc9szacMwc9gAnspakywfiy8fI/dxqgiNIld1DCQ7irLNWn6hAHiAYS3ZocW//pTl+
048750kMOEHNDG9DYKcJATYxA3RR5s2RqFer1AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
fJLMFqIZfVPsSmGW6zC3Xry53Cu9/EjG+a1OHO8aYnjflfu/yBfTS2ilbleEYzHMN2v4hRCEZhrp
W4hX8NgVPQ==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
g0ZG7kwAqV1vgoTLBhurLaT4dybBIxnawe7C0ePiTDfrImbHjeYVgARriMAhTmjQ8uNFTiQk8fgI
8deVo81+FUg3E/FVn65Mabt4J5k8Gc0OeViQcBH2xXU2ZlJK1WRwqgE+xqvMcYEZy+U2ZrptrdPF
/NP/hfapN3ZtBXfH1wpNaSsSaZvsNNqOcbgP6wdDBNIxFuQ7QYKVIwXJTf4JhnWQEu99YncDcU/Y
kzal2Ip7MJ2XrUK+ltChvNSXijvpGE2Y3ZvpClhOeItfRYOycmAhnSr3zc/DenKY8xLTb3d5oHeK
OBzO+jX5/+B1d+kRrz0Y3DbqCTmDcVUnC1MBAw==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
BOu5W37K+fK1maH7Ms6vyNwtjlfo6nWC0lRtgGs38pejv4ZIa6SPemcom88bbtTI92vlDYH2u33Y
UJwhcGpXot7wcEbLymquAZhRph58YUAmSBO+ffAfCLZraXvVNLdc9/4T9KbGI7yHNssf3ErvswFU
V14fKs2s1d9xdNcOfBM4y0KnLDTRh7uDfo+8jATlv5jswFWS7i6jivMiB6nPF+dzvaAFOiyykPUH
gN5QBsLVrYHoi1NKnqxek8+urm1Zer8RnoHYiG0EroXiC/u1pI+h0negNDYuLqe9RWg35G9GsGLl
ap+A+e7tNrO01zPSuXaGiyhwvvw6Nhef+mtKsA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
e+KDHtmSgioZyF6e8SbilgUI27IyKV9Ta6tb2dqMspj/VssGqn4TMTm85tAQ58NMU7Dn3vex3KRt
h+lRWCdbJCOEE2AkEDG/eylcc0l++2incGnX+2pap0UY1i+US5rmspejGF/1GWW/WqzI3lmIPW+l
iRzzhvDsApD79CerWUs=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
PfhXUTNVbolEudnRydFal+lZm3sw+70xrlDzv5uqUhJmiPf2AhsTduPw/psnp2RwAlQKiLihb/JE
35IEk0tbMn7uXvKkKMbGP/aRvmetSXH1Yaz2A/H59qEZNXsPidqVu/7WyZjSkNqIB6HQp5PqmrGo
rre7OdEEx8shRFxTJCPM/UznNBAbPOya2xX1z34Sd5nN10EusGNRVkkIQ8ij5VIyORQjXUmRnyrh
GwXPOEIfE5RzgDglegQ3QDubiY4mJctW3+7jwxjDv3GOtvD1fFYnj3LHnYlEdCVLWUWsb5gZd/05
BXr5ViO1D4HaB33KIRVCaRNsfnGtcRa6mxgYtg==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A5uLJyFaLFPE7reOjqyD1LCk5KvH/8DUbNDgutJj/47ExH7QEIEPB6QcYJQ8pF/rGE7OFND301e1
qROBMCHPPyv2C5spcdvbufcCIWuvco7CwPRLqjh+OKOMpS9PxDSeMkogrGQXTBZf/UhpkZSJ4I+0
jg3bxfyQyhGUADKK4mQSnqUeW1z6khAbafM6oyu0UOtLNU6MeOI/KIq9b/XZKAw0r7avxuNsZfva
F5yCbhgY6cPOVTmlbCXyQwClUZXEczKoskEwcclpay7SLWrkm1+aifsAHNW9gd/ScxAmf/i9OZok
QFjSWrcTiHsB/BuanAPVq3eq7iXYsCDTC1vDLA==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
I1zXrjzUy2VrbpzIoRpP6sBjtSbZt+yX8euQcG7mq1QEAd+UYdyGeE83TfWQ94MoM/FYrnoEcX/y
2IfP+yvSiZ87pinsNlakShJDAHdNxDVLRBEwot2dBWNTgoms29iOODu3g+Zv2i7m6UEKkgWORwdq
WvFlv26N2CXxs413pcY=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ThRLA5434SkpFRnZxltp9SvmijNC7cZS4edJ2r4ufzeHzD/X98s4BweBD4HY98Afj7Rb34KiKPQ0
7Pu6sVPr2AA9kXgC/kI5QIidbj8vcZrdCYmggiJuynQ23h+opYb7zENAopysz23gqrLwIfT4rtCP
hcb+LcCMJxS5mkMstAI+VufoX5fI2Vk6gVSMf2g+NKQflts8T6EyTHbx08aXEhhAfuVMY10WXwgx
ot0QHh5QMqIHOjtZCjndXjmL1L4r2jbNZj/kDBS0Yds9miYp/Zw/ZWXdTEf4d23SzUIJMD/XeceN
UnExjNc8A+PWGMyCcT0PdUd3xC6H4wJdqrZodA==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20608)
`pragma protect data_block
u4pcXU8FLmZ0/81Zn3guaioWGbzS4GkpQ/+kyU9jXsIR6Qx75NK1ZzBhsNkpBanFH1DPXl27DJae
IPicwnxAfGYA8Z7oi5jDfSuJ86985A6Iy2OkT8PQJQYGFvdK+yhoIKgUyFKZwbEglinm5pHJUMR8
+j93V0W32+82c1xjY7bAQnubKgx4b6aocKENdMSg6kuyffh8Bj8d2/DSpdYvQRzQkWTBn9BfU0n9
tsswarHOAQ8fZCVBWemXCHAnwFsBYsrcNCJd78bNEFh7kIhJcR1Bve/lOrNC2eNaaz/Cv0fc7xO4
qVyRL1pWLE/uyB5+PFLhYhSPe/u3ZEKshKHoZQv+X6oao7y71eZcFP8b3mLcAUhIwOTnkPLtwzIl
HWzLZdGQ/5k0KazPKSx3LbOYgiHIa71I2a0c0iF1zjL3PXVuVG9ChuDDazJpYJBnzp+MCn9o4AbY
+UGryP5bjQzxBg4ZsnThAHKeVAAWNp7s55xmIQy0jehA/tVb4+KdhSX7phHW7AtBae18zVXoG0Hs
sp6hE9D7N1rK/QVETueVVUY7AZxTDhac5wfGGjO2l6iymBOyfhjwEbJVNzOQUS0YEwk9dUN85bho
hoF1weUMAe1HIkXXwk6DxA76YwMks0ZW505/R/jNVv5d/nZjg0tMa7jDsEdtLWcUkkNyUoMePT+y
htut93F+Hbc/o6j6zrgfI2t9Rrl0ZkNvDjaWOfkKNkofVdq0l7/XbMQcxr3zc+8dwlKHCZksYvpW
GI11erCWHDr2OBkOU9KpNOCuKHHfCRee/l4l86M223l7ZdG0Fv7QkTpVQ0H5WcdB3Xa870msYn1G
udXyJIGviQPXxfHeGbGFqmnEzLj0lxfIQPba5DCUOiQspOeudv4PBlUAiiAgfTrt9indptz3ae9A
iLC88Cj+kshCv5uD/9ak+bk8uqK6RJlXZPed3irGZxbv+4LOaixx2JRmXoahStA1FOf+f1uezyhK
Tma7W1m6uXREw2LBkGKrAMWvhPtz6uXPyxErBKXPGKNkc+Klf8mY0hkCjSMnibcw83gtxEaT2fJE
+NAO6TKQF1KIBLqbqI9FcRRbRe1iNFCjVzlrSD70VUQn+wtJPxct+gHsGzUFlPPvFZuebpRlzJNW
bcIETwQqM5KNQJHsBli5NanyACaBYN7YMGgDjUjQpDY2BoRndVS+RZcPuS6xIjQA6NM9Wrk0ASuk
UfNJoS7/b7j+k6JOcT96H1vmJ2BcW7EsRxVAAFbmDAwDNJ7Nsk0aUcXlrLg/eFI/IhMAD6sYkjtB
1RnJ6am2izsH20HYMOeNBTDzr38izvo/xVEs7YkNcuRdtsRB4dNaGVUHXNoDVbAv7zkPoCcmCSBc
iRpeQ64nqx7zFiCAHpE0x3+H99AX6Ua2RFy5wLCuTixF9IBAEVeaYfAekuqUoXefXL+bX/FFgioK
Nh5WBAhCf2RQBRL03shBClcVnX04Sp4+W5CiQHDbpkzuG2ih64tLlm8QKNEguowvazN9VNhV2elx
hjGnSMHbCyTAJD+DrrODHdv6WVlF0SeWWl4UVXh3MA5dOITo/7SGDTA2qd37B/5DANZXMdZlKYgp
TbiyuiaaHqQFuGi8pY/8ImLx2bBmtnxNQJse1VTGDl9Z59WHy24FAJ3NiJhHD7WGgBXk8nv8xhHy
HV2qHgscZu5+NwAHjWeOfuIJRhfYNTrUtIDa7BMts2CZEzbLy5WwznzbkDsE8LRPDXbJdmtO97ta
Ofw/JATH7kea8J3owHJ9tHXHaM8IsqZP7ZBzC3gLVx8YIsAu6Hfw5Gmm6SD9B0eM67UxWVVMJYGx
O0UKUscdi0ZBpepZw4Vm7EL1U3ijxKqistDGvIfcbrpqPLE7YXvRY4NMoc2gPaUQDSJtVMWal+VF
cC6NFHRUHp9zviFmfskB/4IJ7VApnNnmH3WwtxXJAVB9i2haZ0dXQFxtchpY4Sx57qnvaJvIuHZl
p1suDWOAPoLBdytVzEtLK9JrY9Ene5GFD3hhSDMoq4O+YPx/1XG6FBtRDPLcHE6OLaYBWjf8x4ou
XFV3Wf9WpX59B1K9ZP5MEmpXkesDxwY2eG5wXc9YWr3InzIG8nNwOSQsu2S9XvbZzTNNGaCqOfFV
M2akmVmKTxGX6zTIYbVti6xS/3/r9i8+VEAoHWPElI1wQZwZ0o4pk+zGL0L2PiHWNm6V7SQCyL62
GtkiAxve20XNtLrXy9cThoFVD1NFXIuKJH2cMIlEMijmvF66b/ZiC9fGZEnPW6NBm+KFrsfcyCpP
JDtbPUhRP43UnZVZM2KceUSsNXQBlvABuSh4Xwp4kM2cBmYC3PMjlRyyXiajzfyTrD78y8jZiEPa
WBEhpdyAgSA+kuSwuMUKiQKbkjcdQhIdf3wG76yjftPU1bAjooYFvlmYwMrHBzutsczK+SoFCyje
30bEMTICmE15lWe0bc/FLkGvZ4R9U7wgy2LP80jiC9DIBUAXmTzPr3MmDXUx+FRwQo5eNyMv8EFJ
ygN8oiRuQ0jdGVXybhelzgQfO1lzkHQSeeb2cqR3W79exEbrV1O02MeEBTre+7s7wfoXS8FpoXL0
M5IIla0JoaN2QMB4N1RzxEQleNqA4JFD9B2lCGXWewrUaRlDP+P76hzvBNF6FspX7kaP8ggCiUYX
w6aXH9mG17h1Sh6i62UUyQmbQB7laYlJ0D/5a8M+enKzx+n3hWFc2aTcRf/DxeRFelOHaTiXSXPO
0b7dt4tCUrUB4GHsd7hpTwxGm8BaBlH5+pyCTMsAB8i8DSzDF83lOfqCKfJARvr2k8LJ8t+3ACIb
xkX1X/fqwoJbtGJur54Hyne/FQsspP4tU1ed/EwFYwD84tPNkywANzgqGS9cOztw6fqiDQuUtbmx
uTWyeqC43dQ5oCFG4ZrIPCTmiLJ2/Lfdzm0EYJweD7n+p/Lw4C/ZURD0gdknYDm7IKb4KXjwLvqH
pIbY7xJ5MRTUtuV7Fr64yr5JJX6E+nLok7J9AMw5UC7J89k4E/1CsQMqtZKN5clDeFNCTkJEZLWi
TYZaa/fuIy2OsoYhI7gD0TlBSSbkpnG1dz8QV59ogSTvdWDcRa9xnXoC6u5Qfw5d8PpE5NWYt+UX
bTpFJ76lQ0cIkdw81BqyVvUTTzGuAMibKHrB0KDiC1SE1RFFVSvrCpriWOgp2Y3XaGD+pW5qdS1o
d47pLMV1qsolr+CsLhKFVXSSq6fFJ5HiY6WjHzmy3g15fYgLdsxGdqHuntYnuyxPrGqbmaECcA/X
IN3dWt7646NCXyJoPRBFFFdkmvRX84FvV9fNh9ZEzWfUD9aVXRuNlNhWsSGP9y0jWHSt4NVlVqMy
0PsDyLJyYSmB93feT5AgnzZaEOyVcFm6NDjYzoi2VTl7enzGqjiwoNCMY8UGoLM5/IhjNwaGVd/E
OchQScHpeQN0toC6daVIcWhk9tovUuBVhMR0nw9jnwksNrUrflxATA+8rH+dltjtzdHa5HuWZu12
5+jUDjVb8KfyEt26dvYrvFVdmXlP5zFF64pNrE7k3WiA/M/r8hyh6DMuiy5uxQFUgsYs95Cb5z05
nlcUdcBFLErjpgZ5NqU7MyVBnE0oZCASBaBMsWghddeMyL6qiaCRAETUIgOg3tu+kcMxF9Olhr3E
kwkjdsNn+dlZaBNmhJV59ebmVh9ys98pa+24/WKIohCFAnHqaDTjF9I1jB+5HO9Kw1idLWqoTUmw
vzTJ/wmNwdqCMxlzkEO7lBxIZwN6/NCDTrf84ilNol/UHzoe8YU5XAJu4OHbiECDuBl68FqYlBev
OMnzgFjqYUhSO9aESd6XI6F+qpmvBqq1bBNytC4vJ/sbQpLikfqq8h9USXTSbhgdW3TIDupwABej
LIZxdonP92bMKwe+7VvVREx2Hf+HMIz4EVs08Qqo4r9CoT01IKJECmq5Yeoqmhkx8Dr1tTGgMfdI
W09MZxv8ENep2/fos2lPKt7mniyh1NiKypL/BS6zqG5zYNuxvnhAVjyQW4jgAyqbY17W5SuXgbN2
nAsgHDOznPjEUYP2ZxV5oCy95SEyTD3/xbr2RR7MMAhpBW6Lf1u8MkVCYmNmvACNSWobwnYwmoZf
ZDCg6sl3aE6r07lgOrrGCCu459JpYObN8NkjgtwN07OE9w7yZASsgY2bUUt0mxienpa/ek0AWgil
lHr7nasjDIHHhaCH0fMFkSdfaqpaKHymNvZmgJyNO6fQ72pHqE0IOFXydAvMsAtBcPGQyacTdiE6
bEIbiCaWtfeal/1zalVW04WLZ32s5Lai5AsoRdaxatXX+wephJOAcjAqQxwc50p9QGf9xTquvCGe
SOqL2+7ONmboANApzv4oAFSD+FBK4mzWPi7nQsye3G0hSAPjRiw+41ABqsCR8H8Rq6dXze6LTBs9
c5x35152pMzsGG8O/5jkFrxsYv0q92z7zthhkXvIjYTttH52XhyfpAdEd/ZPW7hoq5Ddjd2i0WjC
mTiZ025vsdOnQiAA/igqIR8Ae6gPU94SmhQYhW2IdldZf0fbv+50NuobbiVi8Dx+FcYBerxlEQno
LmK/VgsAvaTrmiezTjUQ8msIqRxFi+V7p8+vFAgKAOmOAbGUapUSz9V94Gb+Zaa8EqYqfrtyZhlJ
jMQPjqfu1rjGjjYkAim/c5XZJZmwxyE1vqiaSo6zZ8JWF6qDvRWUQCMbOeq/LZwIJwMbea4eyZGa
mlW7gU2h+yATHB8DMfU1dd6AC0LvPpjNYC8AG/byuR2NY3DlFGRtzHngi3hwhIgYqQ+Tx4RP3wUF
qauPUjDMvsaD5F0vXZmjAxdHit2rmYlLxmgHvILSCpQJXWMIgM+6Td0tbec25JV18HYPGrZB5yIr
/kb55Bs1qXeXGsk9DjaRec+leGQFzB2emRk5fz/WguvrUe+P++CHoAyjMwP+WDjwtnvuqx54W+3j
Iqm2cjr2XpL85Dih2V38MquIoTktxsWe2gx+Tql6KlmTNyYfpjfYOUYRkVVYHe/6gPjwNQisPHS3
rOR6wjrd8Pq4+3nrIsQvTpFstQtMQbC8Q1t4xK54/K5BWv77JP5xYgniKK3fQl+fQR9OZhgv1qEV
4rpcRr3v+2eqwoxPGKzy5+gDaSSmPMwPn0lgOfpAfy0G0HpDcnSbjqjy1hoteC4jE93oDvwxPjKm
82xa0dzXTRM0/45CinEeDimFUqNuCdKDPxyvRtMujxtfi8KY3pT+nltcuVt+YxQjOwN7UmsO08ML
kyr53x+L35GQDMJEtE0Upmv7y5QElW9vN+60miadAseU9nBIGM5FKgLIPBzaTC96LDHf+5pRjdds
+2feuwP8QtBlo+VhL/zlZ+hzTXXIy1FADAFkl2p2fZ2/20rlqrAzjl48ADMK4E0sSbZ8u7m+0u8a
cTefx1uzf1NVbwA9fGTvYD7Oq2ornwFzAxhBgx5qH2984ZKw2jZDYrlnwa7la7NfBLTl5wu7/17F
GvCKQ78Ui4yjneSijOYCTJbShz6ZPdcxFIr/s85ww65QPNDRUtsh+DFfxXnpGIvOJAVm0yyzf22b
LMWu2nyObvGUNvVxyRKUOZ0KqHu6SLVenEcyC+uuyTInKRYcudxyL7vv44mQXmuWnwpYM5Zrqi/2
eqnOpyNrm2Y8F1pVESomSWC6+r4rOZRvyH45nQHAt7yr1tSKs2GosFrqYMALO7KuAiPEcN/UYcOy
Wv0X5oHuyZjqaDfBxYRyar8IQSrakRxVxalQRjQH2Luqt/ad2Uz4TBovLdXUJrLCPbqeThFmuI9C
favAM/dfHBETe5yxV2INvUPuT2UnKj5bFyVlI1pPMqeXIUI+KjkoMBCVFqSn5N87TAC7M+VC6dI1
Zulu9A3RP0V2oB1mdVFrV7NkmpZjJye04A1saiE0onFMUDbFVZJH7SaLgZHt81ME973ArToJZOEo
MKLPEFqigfDqKebWCu9kUb1/R97Cx6aRw0ereVjuxpgYOlQS3aDRyY56c+7Duuws0mNq2qgLJwRV
0AA9jBjifcfXTMNy28MvzEC2i7vvhItSypwFodfVW1sYSzKF355sgf0/VwS4+Xvhy8ezJxGkkLIU
8EWlcJrYeDPdu671Bny3Fbk9oY1W8UMgYfMpMwo7kPrADRLpX9Ml4JOb4jpQNhljC9xmdkTihHIo
mzLXv3G33eXuxKNVpGnafAZ05n+R9HfT9SYesBbOdNBNprk6WeI3dTYVofYw5mD6Wh1AeEMB0+qv
SkEjzjsN1ZPAmGngVCl9HiP6Ys9o2iwOLdVXZxocT3SDG0YsLlKaNR08KePsxEhPbekbQoP3P0wS
oBeNfRvITLdIKLgYPx3XXqPgCobSAvqQwUU1UQJ/uM5rDYuwQSNFK45jidXHnu9jOUl8u242nuwQ
A0BO1OEveqg2/iCGlzR1VpVoB5VLPZCwWYqLnLz5kN/CPdJUcHnKtElC1TwvljwMwKLmear0jSA2
5r+tP3A3wWYf2WiZKP+f0M/Zu7kYqyzJmS38LmhaB5yyxnfHh8nPZa/BdnZFa14/dNHCvVvEFBQu
muCOZuCwM911aadAIrmQB7zXp0xEUrA4aFEEOCxi3taMS0abu46Z+PO38/d6BHJtVHB0qCOqSF9A
oX5OEkdCt5UFtwukNfmH7YjTp7S/sVIh7Ha0jfWkOdBk21U49wp9A5m0CfeJGXTNwpPeP1XQlJvm
vj2hc8UE/Nb8rZbq823WgfwK53GG0LeSBRk/F6rShLruBFntFmNe0Dp/3znD8xIGbsLHZ44zMJT1
m4d8yk2TcnFj4IODA6VS5pekHbUyxwg17xQwrqCSOQBKRnhN8eKKHxizhwLvZrEpLA8q/0cgfTxd
n7N+f3uOMvKRFAD/7fwR3g23CcsJRUZ26cNzZjbA0MNj+1bz6YG979VfNgTS9tfcsMuzCeIfMX5Z
OqkpzUdp9kqf+V7Qw2n8fUgSrGO2/OgsvuJ/pVGOCbpDUUrm91ip7Z9e1EcIFyN8igSqucBMktFI
h7X1LvsPgj0oQ2rFJOxxx+QsixJh5Mtp2Y5cHwJldj6Mic7B5wuLlARQTEp3P00RBFDo0/HOv4rm
8BsNmmQg+JzM0eYLc5v70vGl+Uwu/BoxzKo5K3dV3/Z90lLJi4ayLrz1xGTRXXba9Wix+bbHgiqM
x5x9haVfZE9RZ/KFFkbhS1/7l6XoqSPzkZWqWjRvRxUZVjHJtIbpQefUvpvFh5wc5oSIaMgxdz9c
cTZkLOSBU2kgl/j1GUPh+h7sohwGM/KV+njt+BaW9/2pQrG9nvhAm9+lM5lRKGRLAwPpKnI6svx8
GfD68R0hhk+F6cEe1rNFYKEr6y4GZSTOrdzxyZSyOP5spTto9HtqHZOJ1FLuVwVkIhaAI4cmwqtJ
gQwTgI/EUAfUyf2hrFn9yLimDZVOMwndhnsTovOZucXj2yD6u8QEhNxjN1JYFxYCa9zRB9vUDUAw
qQLwj3GnmpR8dE6C9vTOb51aHh4AQArKbSJNjBZVt6tLMtyNeE2fs75kyUGhBCTNHAhocWhAF0yZ
lGIzZI9JVhr5/WyJ7TknjR5C9LuenzLcH+iaZkvA6xH9rKFhLXEdO5N/smqKbuGz75093B/LQ2d8
9cQJt/BRKLuEm7KzHjbsg2E9W9Qio+H64vnbxipTJ3GTfEzynU1wMr6T5PQyqM1969bSxLu1WplH
6yna6cuGQykyHqY0YBaagF8zprFiGIrj6qfvW5H5dVu1DpZ1lL+qJ4rUnsemAp7+AtxhsQpKmDJn
aZVWtuIOaOegpxaoqGihfZzyJnVb5qKd3YR8W7MmCjTI3q0R9ZjGlHYuA1k7OvGvHNIrcHCmrcNW
apiGZ0xnA0lNFthR8VlTktmvtW8wMtMGLBkPFu6hBo7OVUoHewnwvEMZCkZg5WTVwpL8zDqb8Zyo
hO8DBho2DrKGZSJyoE+1yZ9Xb/tDFmxrq1SyQe/4uzVdW1DrSWESC8Zn1lJAN2W6l0lVknfTDpgk
Hwu4h0RCOyAMAIm2XJnxIvolGQgaM3AwJ+elT9lecm3VnnYwcMQdluKJ8DeKfFqYGc0iOlhIERLK
4KImGMrUhqvYYtOa2Up/1uuV6MJ20WvAD7aRoaV8CfmwTCdIP5Z3j4DGmEmWKljD/Op/7Pii4YQ0
HHKmq54PPJbww9SZcHPSn9xXIZCGbu76TJejmAgvnVKBdY4TCoAI8vPYt58Nabyd92zJSIYXeLrU
j1JoKXQJals73jIv5NkOZJkjAJEtikqHwOB7tb2LaMDHVtJurM6vxbPLotoEtxfHoW8MlxONGhfP
AGfk5lGvSDEApAQQDbTZflYyfMPZx4VNxcUmC080PbnegY/IbedLPVVObvXRvCljGZL5xSC+Rpkd
zyDh3i79tcs17kej4dXpeAGrX4/6LC0YSRcuEwh6TAvZLwEx+1HMnUFSiikV4/B4gFfU2XE6Iifg
dCsv6zBgqSn4YL4CQ6dCcl/HEAs3Q30sb2C9bhGerxO5/Xydz+OJNMXZyrbLVaJdLYStQuOJFMBq
8d54zV7OzzZX8MZOvbr/5zdDOsWbEO3zISZKHFi0v4o4lEJe6o7deyKqqQK5wxAQxBjyU8s1tHvx
HgrZe2xUHXN7a3pmZya86ni0iGxOaXVFMlifXm5bNv2iP3gCRSLP5UrpAbdapwiH4cawKkPr6GX3
QNPq1DRtoj71H0rcrk6erQ9bvwm6EYI+ZM8b9+63XIfjVXRuI9rN5GUHhc/hmKtOK2XSKJOUwqlf
h+/O+GRvMOdKSLINc/HYbL6ViWOshRAryNuuzG2fJBD2jGR7Ns/KUAWmVhKIxTlsiME9afxmHFZw
HCfbVaiB7DuEJqhlwkr7jfdlx0eZUChVPAJ54q/Uez4zcdvlpnvELzP32Bk7DfCoo22Y2vOzy6Bu
oaCoW6AkG7wGFP7ZSiXo0/CSNOW7DGKaZLBdNFp5K27LD5PRy2aTBcikc68C1/ela55GyZDPBaql
3cStY64HWrD7aIwUwatdT+haXyThk9DDyBjJRxhRyj4DgrbddPWeuxbfxqc4OgRKgb5HH4NxjPpV
NXqUrqUCnWIJet19ZBFzRbCDTAlIHdXe18QF2Kzyb6xhz2pl/AROWL+hSTbIJC6vYyDHfaLZ5VOe
w5eoqnd5XnGK/kcENwMUOpXgA+65QwXFR/tRM/5w/ZEhUsdoYtclQTgZzNqc8AenYNc7VqhNBcdz
JrN76OLFMFF/Ww+x5vgIdZz4deCo9ru3Ro2nAUmXvLEQyC6qZIbmDT61ChY6XOL16Zi9tATcD/Oi
eBeGX9cF/4k9EJ4ZTheUvITzfMO/3pYHzW2FKzGxRaP3mVBo9A7rCqUjFO46vp9AQsuBUFx66osw
FCneidtD4fTOK4NLM9p+qT+9qUMBjNGHA0kys/6zdApug2IvIyT5SpXTfBDkMtO47pqBCr+rxbym
A/8AL8e/cpCKVqOWMQSxTzI8CW+jvGXdawkaykllSdX04AyNS70A0XfBJwl3Z0ulo8lZVBC6NndB
YirWQ7PhoPZ/tHkUX5UE4Rg9UtA0uDjogXr9GDo2YkKgF/EYwQMcdF6H0voFdbC5SUZwwHDzwJtA
yHiJU5JG/sMe/R1WqZ0oKu2O+7Ml7i/4XkHGnjFPNDv3iRgZLB8bisDipzpDwor8GAp4SzN+bl/O
7pJZmIlJttc0FItX1JRAlvQ9a+z8cBpLCDhDUu5y0qb9fzQJSLCGc8osphoy0pE5QeYLhqd++UhZ
qHUP1xPg8zE7UhEBfbjZDjHClmw3KoQyraHzSpEifRPMpPKu+O/tBLGoTr0L/O+Do+VuU95cHKb0
LfdRpNDb4zMLeWGKICgSCX51yLeZudaOpi0p5GYhEpdo8woWeDrwu+MCjujdS9JsHhum00W/1d2p
rFUcxd2f0wDVWMwBjXbzy0IVoP/NP9tsJpRVgi7C9+Mp7X5SP3K4ZM9E5sySets9m817NHs//bi+
TFoa613L94BO6jGd/KTIGd2volEIVbqAAx7KO+nVwp4npUtyc9sJ2iZDreryu96U2AqGPqaXI3g7
aEd7rfr1U8PI4ngar3OKgX5Mt2Id25BksZOfrtd/WWb8lkq0K3YlBLSIxBBr4YWAXe6Ztj+oZBbp
ts1SCFiAzi2IrF908fyxhKTuLr5AiJPFf7w9ABbRwmnPDq50zHN4jzD32fhf5uoZaKgoshWKbI3O
/wcsjG7226ZQY5tQd9rZvAnz1Kf5JBqy+9Zm4YP4xhhu0X04qi8BxVbs2X5LQP1qJmCbmI3E8M+p
G+2XLoGwDiTfn/HL9gBCzfDfpffLf2EE+LROamM02FoadtnVmAdrgX67MsjU3mBMB608/VROn6og
+z/3wrUxjbzV6X1TyTvdBo4b5khLE+sqCB8c4XVJRqk5kXn9Z+Ykl+OPejR5dHPRlh89Fu/ioQs/
cCiU2UgECEgeowL74tv6bEwejzKF6CqzegcD7Olh9KeAYlwEKQIF7Ll2ThxR4aDF8w6hgwsZ2i7E
q3C5hpExlOtTRg6iWsPYek0rRk67JBNzJKOrBNI2BainW9gWS6BF4GRm8Nu8IGa9wULPDV7ld6K0
0jWfJlFYbSzQk3VuetdH82k0HsrrKZACl3yKZYqLo9aGLCWGwS0oGGG2+S24M2Kfe00TNzJiqLnb
mQVGk/iACoxHukp6ghPsGSO9U/nmnD4Ht0E/3g+sknhR+Jj0npqJ1JdGCBxSTrnhgLpFzWuX3swg
YyAfqHAJBHi0ek2gadBIziFh1Yyzq6ytfWF7FHGN2LPzpExaO5tVdLyR00k8jImwFol3quamA2a/
L6HDtedNs7cr9ilMKab0eSPAS38K0iZvWYiiOOjupR9qhK5frKwVji5HtbyFBffh8O2p9IwTn5xS
gMMc7vtLnEnSnJ223hQiO+vv4OszKwuTzmMpVob5mCJpKRFFn35demA4hXpQ4dIK+JXyXotxac3Q
NazjfiLUJXZ+eHrlF2szB/sxAhImuHftlGmSsAUXPEEH2KgN6hh7YbvThIhrccff2nXz4/HJizGE
FAWbDpsZ/wYhb1NTOPU02W9pk5F0Hg5cD50qbUspGmyWYPuxhL8x5K0lNTe2j/S6HVk8YniRtvqV
A5YCo2ISiIB3Uha+EO4vtcPdi0C4n7yesBtuSKLxINFx59pb+VarlslEW7RK79DzfOUgd3cOfIY8
vXbCHBs/rOuQT0XYb9kDrbC97KSdE3Pr5WhnMNIX+bRMcFlVfs9gUz6oK7y2heHJ3fXKoeyqg5+d
GxRdRB9z70XAeXC/joSDWYGEw+AAVmiPpXcOzz2C0zT20ur+CBTCKm11ynxfPqcIPSqKBFFxmS2N
DXmXD53VvQrL0ybCXtlKC674u7SjCiGp64WrOhx7ZRcATm7h/qTqONznwf6FX/mAjGgl8x+ngnDQ
7EAZTjOTFTM0wrLofyuy3V3Io4UgfbekQXPGamttQl/cE3c8OaERYEsdxYJCzXWGwcUrBwmCgHMV
UCuAe/B+jyRnEEpryzMpRN1xQ28zmWjPql7jPB3IxlmGe73zOOjn1sO9ZbayDJmaYiUnrutyByJe
Uytj9Xa27XsRCjJB2G28T9QLZYwBaPz3quDn6CZC5lpOWBQPQtzsxBdBhfZdfSACxXYWt3ejl+UN
q4KDxIsK5ebZqlUNnKSNVJB+6V/3b1yRug7xbdzmFaoUNtSljk+k1gBGcHj+X8WoqDentlmgDOum
6Kdiu8pKp/yOjDCSOt0JjXD0I4Brwl6MpVUwPJP4txKzBFrmhB5ppiGo5Yag5Djm8WZWehUUoF75
U5gAqThznYx9spmQTXSsCI+vb/FzPQsQqqjPaTVE59MD8kOrpW3ewKY6P/V++gd5lEtkA+ZlnqV4
WwVp8X9OfGzjnOTquJ7hAdg5BJE1IK315pvRHtpBaOywU5NFWa4Ey13Ajxb3np+bwVD+MivSG8xV
QTJPLABzy8XLmxpzcWS8cPTtV/pqMbGTZV9ZBGB9FFabNHW78Fy5W9yvfSk5HiesnURM7xtCzhzA
xHgsIAIWeGdgvH8HTwFCqP40TfWbKYLKFbzR/8thD5aJ2jNyaFdsE4BiXjBVhwztzKMasegTQkGo
9K7qvanbHCjVP30B+12joI50zcUz+hRGNf61Wmd9zXAtDMZxAANJ1GsolmMD7nZrzoeVA1tbEcDO
Lb1iDyPC+ZSTl3VjBrPrbamUW9e8xki5ZqVPCs3OISwWYslml7OtNRKsEBylG1XyosC2A0zzSIJ7
wh11ezqVO7OhBtNo1Cr+B9XSB4m8kTkM3RXqP++iBDByxBQ9VzZqjlSgZptZS9K4Ek5ka7HeOjSJ
c+ol/h1NfUTvjj7mVCnzEpLB8GJLLINZMiV5z7F1ppzlwbblGR0FJYAqJgE6GMlgK/kmWrrQhBBF
C/zJXspQjaFe2MxtZqNydvVk+g0ISKpkeyl2oTXZRVcvfI0SlFklqKq4s2hERWGTXnVs6oOj+eS8
fS39AB2yk4kzGeCPefGaqxO6S/TDJJAed5Q3grdvRq2DaqMhYMsBOiRrwarMibT/RDh9YNc7+mAb
ZstiW70Pm3e7n7q19nLhp1r+16FztgTHyWmVwxwjTUkGrpVWBm/35bs6fO8BUNGpxykjfCybpCCL
Ad/Eyoqfl4xGD3vzY5cGxyq3Ern6q7QDnqgkNCc1FhLRu1sVi7pMakNbucheUP1C8YyJNQNSKZ3I
41hooAyjNMM9kYwL/57QNCVL7rU3G5Yjv5RIQuxgffTKGa0rsdQuW6+mkgnopgFJUAP87ZZmi81J
y9VrQYxNX1xdCQYnijswzaC4TreD+goC3z8vt7bPXfrmzRzTsyHNgRlY2OuQUTRFcpMtSJV+fuCo
1v5yEPK0tJrpdJYmyyhWUA0VFbt6ZLq/GJLycIVOywotIMC8lNHZ4/7p+gJ1kIyzeX3u2tiL1a+t
om/NpwLk4Fn2mCiLcQZOFbyohqeeMEPbmttemC/uq95s92wWn3Bt5WXgcpKXF6dMw21TpANfhj7X
n2gl0/7M/pagc2BHr8NonyYcyOiiBZGoGcJw318AOz9+uQ0W+iW1YC6joCR4UwG5C8hBd6fYFnpL
00UM6zIsnKp409AYJSxi/Q8PLTTBhTkgk31fTK3to+HOYL/vpuCMeZIDFFB4TORhks7+S1DksWCn
kIjRbXZW0sMuFgydjBheXbvr2UsL0qxlE8ETFUS/6ZYpenTkcG2xM8YXCpV9pZYpORnG146hWYhY
lilDPWgY8PEAxRCnmZQqg7HreszvFtGShIW1mRvfy9WcJq+RYRiZ49BIH+ABs18hE+zlqHKiUBAA
GEQr3046sH8Da+9X8hQXKdk3T7gVilW5neTAP3coz2VK55N5GbrcoEbfZI7f4A0s1t74AHLtpSr/
GZTWXy/bn1sBYCIqAqCh3Q0o+Qv1BxB24A5Ez+RRxvXO0te3vepliC1yAPDoheVAe17h9PqIQHQE
wxC397u5wiKDA05irTrlp4c4OHK/jhHULCN7mNFCb/vg61aicNoNi3WwZfmOTkO09ToSQteqhoYR
Bd3lg/LStcctle5FUz/BdGcLbpsRAeCF42odrEbT6Udjey1v0P4n5Rp+pJPO6PTrfAeuvii5hHp8
htXLnp8NGIBUFV41k300TXm7jRpdLncJyErXlEQi5u5FbC4v0IP7wkSLsx7hk/qNTaraZalQZvvh
+x8toEZk1KgPf0hFbPRJuEQGJB4NoHXJm5U12mboX0ZR6Njc6Ot8mZ+0GzVms3O3ZVcmqlV9q2hw
rvXlPIHIIuaemJ7BDG3bxnh6KpwFO/jcfwmoSxKkaic/ET/pPcufO2KZSUc0+SBW/b86+zWQV0+Y
dxel7fC2Vx5EqdYUZkizq/PXpw6S7hZ/0SKquuepri/HP3fjU0rw2VPqKScA6GRIgx350qS3o4J4
4r4Nh8Nvpeu/60NzxKWo8VY/YnBKp4T4N60g+Bo6A+MzHuKdhFyQjVC5Ca5hEjGTnSjHyh/WN+h4
o9STMuNuv6Lk1IRAtIHYL6VgC+Z+jC9SGfYEytmeejYgl/mVoNX12LWyKop1HB1VxEDaWxVjKrL3
QIDEmoeK7AqRAVeLRKbboRO8J8hRI5A2SYQiWJwftmY25iR3v3rAQ8q6G3wTAilzACeQtuGStaVb
zvY90NChh6MdXRDKKHGud4Zc+hJQPvH0vyBjSaoygSYsVzUwXYrFDhWlqozWLfOSk4NU8jqPkWoA
aqahIetfcpB66nkSvOkUPuvNguHW9YqR9cEKKNu1cCz2W9H4PTO1rfxARFM7KjV4UHr07HxgWFJa
H3Bx/6V4GbeHcsFjAQLW6/BFyNAQu34S+Sq7V8og6zdVEmfRkmSVVh0b7uXMLXJCJvYIKxFpLn3B
tm29O2czaBkTqEMHdh627u/VuYwjzLz+Pt1HTh1BGU6ObFfHlES6glZ87CnkkjFBJ5tky5Tr2qLD
kWRXkWgCMA2wN2Q65G890aIjTWaM61s+T+8qTu2pg4aIorSlibgueFvqAfrY8reiVy/dUUWSleRf
dEfvvLqQwXdhXRLUoRfUS77+nX7dx9YegPl4D1PU/WqWkHn3wOMGCRUY4h/yHvR1JQFEmAQkminr
IuKJv0yuSJZLsde2grbYZG4XUYfyhFCcUa4byLRI3H6rN+5uDpgxllbWeCmXkyB3fjNGbYHZowL4
DnwkHKiXC44CkQac5tFFbfxdmJP5B6M85oOB/bS7HYlRzzeZzDXcmluCZOsVt+F9DVHZAhYTYkkt
NVWGVCQUwb68IWpIRHneNS6wUGqpcwDafi3j4ynCRhn+ewt7WoO5bVqhPJtrIFWyycexFzaWuSQA
5YpZjojMU3lffmgMnt3TRxw8vohBPWozNcAJ3GKuOr47xsLEIsFqef7i1fGBT6xZG8lutEJMmceq
YM5HPJEwYiS0dQHz9grgPKX/eBiKgW+9oHhYnTqDu4LaaWJ8TK7iwxrcC/TSfAs5RAi8BPNkimGw
J5WFny6Fw5I7UXI3WhCL5aBvFg0KyxFW1eTp7I+7q1oIs3J9YeOk+Rfjisz8saW6BZ8eZdHx2jlZ
ApsQb0zJcXj/RfQjQheQSyHEP0ORpi/LCw3KcD3dgVM7yZ3y6/XCxIDvXMJ8CvrsCHwSQSn4O0u8
HUBNGnFh2PcormFIQqhF55oTB7+SisP/RWkQNfi+QKqAnm2V0hfadyN97n3O7ARF9Cjd5GIg9Op9
oxNqDW4Xjjy4RMsB9HAb1EHWVtez9cTNIIaW0NyhNd18S4NwsjgLC8IA4Z4Qu2wIzRysoSF+JqLY
E/3Nu+L3D4a0ogNW6KB1l/YfQbFQk12b6KIUNwp6v93OHg2bk8FPqghxCojMNrBDpBjHZgVr3BdL
XECe6JhgBJzFo7X8UiOheLzjQjehDVJBWLWgc4MZnRHBXBylRYG4O8Tv5jhXWWn2Hh87vsiHqqwI
LJSlLi+xcMq6IbFi9Xjp5J/dWf3u+YXpnqJr56xkKEnLY7FGOUEsJ+KDQ3r8x1VgKOXaLLtHF9ZL
wyc2DIlYR4kvaEhF/hpJCl7pjr30cznWIfyNYqfL/RbsbDbyYdiTBd5N6+bXYWmZg6tfA5r+a9Pc
87xQ+pXwDc385tlRvfkK8Xn2Cti1peLqI3LIiuuSiKnBSsYeyD9RzcXayV37CJW8HrjjSBkRr/zo
Fgu9TGDlbkKxdfveGhVLRYrfi0IBmGePXHX7rXCUusROWWtjtALaVejkwStgM/asnOUPt94dTIES
NW/mH0c8gBGFBqZz0APqvjKTMquHR5ETiyTriAmwnMvuIumz7CdFqOXtuzAipuomYRufzjN9C33l
GZNFmeCwoYJbEUhd+stFMVQ2ekwZ/6pDrHWecjMexYhnp4oNfgaePPXZBonqVbkhDxZpmD/MV3vg
BMlAWvxzVIRdT5zcVJ9KZJkXx8xvNpZTKJ5nesnqO4wS8bKXd0d256ndDhc1PH5H9L81dmcu/YwI
AbZdDY4PqUSM5YwQpS73pzidtrA022kEwB9T/E9mrVCNzTLeH3V6qCV9l3VF2AgLR+WhLBzzhttj
3FbBR0jLtVo4ffbJzeui/oA0yZuR+uGqzjs9V5jBU3t6nF23bVnqLUkYJM1XoHDgYqqyrgJ9Ne3T
frzcdojpipF1e33VgOlH8apSggSrPEkRT/h3EPdO6Od5uKbzFKPkka2ZVyx88g4Fbwf14h9VGCiM
3DvMb/xys2W0MIyzX4AqgPM53OCuvXLRB5KodKdiZLSP3/fWnRiJtmu8NbRVVFsJ9yRfXKnMZhVy
I04ZXHE674TIcbIRsePH44Ck5ZAW2iklDXqfaV+MV1fPF6wqZdClr/AExkaTT6eILCyicu4AgaBq
0ov31R+Vk2uaMQVEhcYIVosf9KYlpnHX8dfQFVXKC8Bfn3u406nEKzVrwcy4S6+yVnp46jh49hTa
PMXC5AcqeFW43kLCMYeweibbbg0wmO3nWimqCMWBNaSwid9ejVD3LwkoiHVPtbPwt0xyhAuM15+S
8Wscr4x0hr4RL+yKBtcQkXlpjG2kQFicD3BLv9hajhqpEBuQkx9pQvjA0kLqMso+dtpQe43BRcSB
RWRHEY5xosH1u0wJ8y4gYt+LvL6875IPz2Z57WRwRc33yuvL6eftGnjpT6IDG80ISKE8wr9+oDic
Ndra7lPl7yBRi3WGD/vCvvRekN+RiwDtLth0Oe55eJdHoWAqKhIH3TeQKPjc7oyHmMhIU363i/Sc
Cl5l71sWHVEfYObuYMmd72fwpXkcRkPwgW9pw69d1L0t8VBJlVxucj5lY+rqsgtD02/vu8WS3Z1l
YSAjQd1gQYcTTCHp1SCBREajKvMFaWJe9+ugLfiwNsCza9zZcoEYQDL6MfgPzzk3Pwy8ulkuwxk7
hdH8/vj0b5liNAU7FmUA40uCb9eNO1xCnlvf5bslktgAQ8MOnv9zsDKVQwQTx12TIfWY37bhXRYc
V/ucAM+AWv6Qi4Okf8ooyHnDrv0/JZ70Vc3dqPJIDEXSm969f4F5izBy9raFtC9LN4cKyH0ss7N9
X0EFQCWGSMbvt866Ps8s7ZQyHy1tZ/LYYDDV1Jg963u+/JhDxXb1LUEn6x++iYk3n58UFuV+6udu
4K+r0TDEqgxTslqEmXHvtn34Dzx2WsdTYopZZouhuf2xGw/cECTDB8xaFhqzodvFKsuHy0qYO4LK
JJqGqEXR5liqfthqHtrGg6E24YwztNHw0zDh+utC1pq0CPaOkQj8Y2jXhGwdeiqsK6dGkr7VIy/6
zpqBBU/si+4lc501Ca1xGe1kmBkVUCE7mP4PjUhNOGBrWEn9wtHT7kjaWqPcXL2PpBXkQ3FqW9zM
IStv55ay0GMBzIDnr3+YTfXbWXiFRGMRQXPLMIj9M/j7SPKD7YTb5lRz3Cmr7VPuJKKXSWwlrhzm
BV001PmGhP03Bs7riam591ly1G8XkaxAnQQO+Njxf1eLXT7X05cdBTa1W2UHcr2Rt5/EhIYzCl+R
tilTCskEmSo6atZKbw+gcpOlaqYjSe3Q3Fhvs7Ejl4FXteGhReMOjAvWNZOhZlhy6fTpaAXsxzyT
ZmVtbrAezqbSMuHMGnzCZzmzGh+S4eIZQ9w7HuG00ygp0p/FcoI1LiBO3fh7G3ocQPU2vHIMS273
c4dj5ViaaYOBQyu6o/CMX3Xy27ej1t564xYlx4Y0+jOCnFEgdL6SL5BkJf3ZK7WtkRc8wirQnvYb
R/MY9SuKyTL0EB/t0WwETAAI2Hg0IJPJ8hFbVlqh4TBBNGUwcpCiU8R2ughPYciObbyAm7W2xiBE
o1XoUEEMYljA+MnUBJkgA3JPqPgK70oNkM3ZIZPZdn2kiDNXCfc4Udfwq9YWoA2An8BFUPWXe3ZZ
x5q3RxBOo7rDGpdBiftbHhngNxCQ0PxBcGjVWK0Q8yAvdG3ogMsSmrhywE1ygZc242UbeeyG7Hwi
/bEhLnZ/R6EXTTe/TH//NTvCce1o0qy4NJtu5o3ArICjnW61a33Mq36IRRMsXZyq4Oo+3AMFxiV4
UYQbUMDzJWNNbVQS3oilGeMEIARruHbIMHRC/0C4+YFw3hT8JD1n0GKS2swsfsyGhjq1pNnxG/IR
mUtZNNoGEAg0HOpntWtM0/w+NvCnkl/ZV/qbe7GiYGuLeVpQdU/GooDcqiw6pyoQditVbboXkgbk
ZkjRutgjNIp+E+zRW236y8T3i3XaYSEK1sihvAmjDIKeYkhJdTcVAGL9RqMTQS86tfrYrhN/MFQa
KkeYYlHTj7uJc4JT2yCkvbph7vI0IyFIkqrlB0q3xAGhkVjI0cwN2vsU1Qn0P85nIHNcbYBZ9yHg
u5VYxmWk33zNJhoYQ8UMEJFqDUGeEFVRv+DJiDn0ZldO7w7ceBFwCLkHWLruLUGzUul4AzBj4yxz
vGcU3C3rwXscNAC+nkfm8z7B/cK8nuOtsy1UAkVw7oPamt86ouGi5LbW2nDZy4w0pv1ZTS+JLp10
m8FklIjuHXDQXoJWpc06OhPV7DHESiIVsnTeKArb0Fegjzu7pElW+W+QU54Tn/JPeP+xQRHyyXKL
P6s7usBcU2K2iN3LzmiJCI22XK2rAekxTQnYZAXYa0Y53DLCaDnsNwfpgmb4k0AzRYZmyafpMucb
x6KLqWuCnxeepAIhvj+VwmRYC5b1QOKAICo8X/67MEwSrblDd2mIAG0kWvnvhPG8mP/3BP0N0aZG
wWAtBPRfQE1F6eM7AIBYTlThc4PLv7eZufn8Iv8YmQOKa0lxnem9HzGJJvjaqFd3hGUJQyiSTDVu
+DaZ+W4DETpOaJOoKpaahF82cwxYuIO2KhhoTZxHAzoOMs2iv+5Rhf4nWLoX5F1Vh2kK5+sWYU1/
N8WmOXCxBpZS1jE3MPo/UPZo1RLpiDs9jiuTq0BhGvuFHKX3RB0dv9HHGyvbRVbVLL1u+CmiEXCM
YxekqFmfB10bzDSNyCSzyG/OhsTkiSzw9QLVUDbAyL1LKMgBFZzqeMmAqyDNAcLTgTAVUiq/5/sa
z2h/C3S5Z4lgLoHZB+NC8DSVaHZpgrXbgCGCvtjz+G2W3sugWVfZQisvW/aFcCAmdB0ivy9c+t6V
kBij3415KFqY0tccCTHilIp/9O9F1QLTzPo8ducnnQ0lV162f6tF2kA8EYS3EQ28MdkNFM0qrnNW
F3/JCx0eyakDSTQ0ZzViW4FddfBb44bW43forT1UoTByDTNlUn9Y6iuinowI2Qqpk0/nsG7i0Imk
zG6xh5yQuweqo11qwy/inM2b8Cp6sotysXADRUs4EYNgtx7O9Avr62cDSIRIKhUR8Fn9vvYYGgoE
kKJa09ARz9iipoIv3Hmaq2+Yvc4eYFS6ZNTqYzDZ+WLZ60+Gv/IQD3RyrFwvjuyLnSLuu+MZ58l3
YQpRg2//86bKgt6+GxYORjdt3hlPPVWkzojV28fFWP8ag4qSF41Zghp5w2OdJGFMZd3+KMCnVmCE
5BBexjpT11MLDZ526bTfrGjLkXfW+ExbNfjOq91A7lJjOJ3LkzOBLIBWEBLM3X4zHu51AAuMTrxx
637tcapC5/RiDNHj2JtVBDaPsToJRwv99fWERdQWQDeJcmNkjoUveYwXjCtAmTBMx/HWj/gR2zIV
f/j9bj68rCjoyJR3Js2vNN0FzA2KOpj8Pn10xjoWCN+G2uak5EZPaQ3g2ntjCplLHbfu9Dn+ydVx
O+h2n+75ZvgxWtb6ml3gWWwOtL+fXJQXaWxT4NijbR7jY13DDXjQbID6PE229Y2FoSMbhzakruQe
Z0HZGceB5Y0Y29JwnxwW/lcsumlNYZfiizoZ9pQ17QRXI/8o/KA/CVvtmnAhqAyBgvJRkqkBG7W+
eIHeVbmt3r/b+Utd2qgi7uZv7DFzTkt8InBJY4z1wTOmBPRj1DRSr/EvA2xUX5g3MHNId2iII/CN
6rrJYf0hGAp4IDWT5KYmWFOaIMQvVpFu9YnfxV3NdwEqBtQCadWndGZWnBUICjozLwByMB/We+Dp
rx4+3GklLu6KFSC9E/YcFfUmATgltZDoh2d4ofcaEgnpx2mVKDRkiUJoCimObSQTffNJv7pgbhFk
atu2OUFb2phVoQLzJ2X+gOl2SKGLScbGnkc+eshMpcnxlswQUI/pQq+ttyGsNWCADxQQ4cBshHCV
/st+l9v2SNM3PBsJAREpFF8iv/Fm25HUrO/nKtRqet64Tbx3GsE9eD/3dyGyAvCMZ5dGOYtPH/vt
N4uyhklDyZqMz+Remu+NXAkr4n1TQoVDGmhehMIRMHPRdtGn+v94+kiYF1EQx9ALO2agaS7FQANT
Kz4Qu/tzpjS/uh4ykPnQgqy93kd78H3Ko79OlqlvOTprbCaySrSd0Pa84g3LQPvWl9WrDldDOBXb
PGu5pxlMu7aF1w/yApSchXDJkZwNiuZv/k+D3H5x9CY0T7aY/DZsjqOQ8O6g36nAuMGvcg8h+SyC
sZd9W3XxYW1pob490kAz2srAV7LqOSCWNZa0wGa7w7rO/dAq2msXAmwLqjjoDlNhf10GNUwasMds
WdGa1xiOqVcoC/DXJ0352h9D58Fn6Y0iv0ThLzm+XWvL3kxUs0LU2lAg8njOPvtebSOLhR8OYgl5
YTsEA3CQxCmwu4Clhh3ahk8AljLwQTJNfTXlwhEJARjGjyUDgto8VMXn+UdIKfKfFTAXx8dCAJGE
pu0JgiJQUvghRafgLve1+SU22Hqmt3xc5lY4IyeeZ8Masn/Kk8J0BfU7uSTYcbhczDMVnHnaC07C
tko/ZHsTCDxMeB/pugkCYFvrfq8kq4Wz9pokQQ2q8ZIIeHCsNJAV3TKm2hv5z6Y9+lo8r8URpSs4
WqI8S1vrratcY7LYGDszALCLzoldCODfwTz/Bfz34hmEkf+vuOEEeNET22M2Av54An57kEp/sQNu
AiNdo0wipMabUYLad5AM3yHybiqaf+YYGjlfdxZkLmWuyGnusXMEK76OEi4R5M6rzqxW5DaRZv0X
V0voXeY/NupV3kvAfGw/UL25hJGHxjV/W4YSvGdYwVetL+daWKoUrCDjP6klZv6pv5sYVG7dkL7i
emjG4C5ldHoT7cEkHYN21/aQI12OLVi7LIJMXXkdmejfCLwIAAlwBKhRDE5BGFnQPdHLgQ0NEmXv
AbYbTJ70uSyMSj8gflkap3bQXJulNIRyjUtlp1U3tkH241vcr+7aahSApICfBLV51N2gRk7paNPm
UHpKbTgiIMU8ijlYIJAc2wR6vWRKWLYfHkoHvDCXoufBb2gg5wZdcNiVSXk9f9Mz+SgATUza5Nya
Ey+VjQ9WF7m3lHbL522OchA2HxMqD70WWoMCXp8AvpeLqxmg2k0BOgTKRN2gdKx8qZC5f/z0lfm/
EgfCltLK5Nre8RLZTKfKdk2DS7j6wRkDreqJGTZ3eJ+AO89oX3A+P6mpxDOE4hHiV+0u0ID/ua4e
RgYyJpzXawgGBHly3XnRAngKxiB/MvkmPHv7l8ZCxXIkZ47wP3GNarGg0sOQv70cmxnP82WTRd9c
6+TN0wOwGFoj7p/b+80eO9sDGAf0QucQZWJ/LRTtB/m+xSsobXLN9Xua/cSqRSNPJvIR5ptEOyXi
kpnfKovkd7EwVeCpusnpWsurcxJ2/sJFOVfWwDldkr4ejmHy8DReuWxBs7FidvOVT9lZwDWDzX2G
4bU9GjL3TmGYbvrREhuecVw/DG777Pm0mbUuUp53HIPpqVFJspkqtLmBXlzCzQCM6vnF6GLsLudb
JQVysYwjUXKMns0tjuBaPJoN7XjhzYrQPgjBLJYLAdfn4alAh5tNBLfjOx7IgORfZc7po3aDZbXB
5ooxKAuHsFSOeAzmKdTmtknYaTy3i+oMbitJcoj7+pLGPH64k6njijGmqvXzuIxqZnT7kcOb4dX1
ONZsxosNVXy6cVI1TmsemA+Rp172ckIzKxAqQob1hZDkF61XvM3F5E3f2X1n2hPaBxSAFEAhZvEY
oGEpD/0GAbEpZBtOLiKVtn6JV15Yz2TVaWvMD40gYjlPvTLrssk8GBLDHON3HoDD99e1kUa9irX5
MBLxyOxQZR7m1hcvtNYz3A4OeHMVGPNMfvWd8nitg1XnQkTcgPl7/t/2sUy0BV2la+SXOlFjzlnM
0S/hWi8D+wYb+JZgMXvI7GDAJYvKZO9CwmxVSyr9qjNthFaHmQVXUc6V1DITEawYrrfwbbAN4ChM
Ri33adAto1sUWlGlBpd10So0QDXx8vvgwduahAiU9N29DjJDc9poEop48M5ErUJHQ3dsnVPro040
h1Wd02y8C9fvCG6ktyVIiufkH9qljCDgdt8sn3pka4LvJpRVxhA6tdv1cYqm2ktW4Y2TEFNvmvGG
ngQh1R4kC1x6VpXPiiGRhnpV4rXFSNN5C980QjEu2vtrP5BxNEq2U89DpwsTnN7zr67I+8UVovLk
P5Y8TUO5fk+Df0pbuTH1VjEVC9lzQvgp3jGj6dbiA+o+Rug5h5cRbEx0ZplfdVImfekG/mrTyOFk
hhmI5jsbwE+3Zpi6VUwuaah1Hj3K5/HNGJpnWEYejpFgyZ0t5BwEGVvlk5alS+p2or3+ABsIN4eA
UfQov2rbBG109NAvdMhNBQl+tFnaDvXHpogCh9IIAtD5ScI9EJwiNZgwBh+Bgz3lUcSfY9j/J915
9KzsGcd++D+pS6j0ks10xoch235QzwVAxXSTtF0wJnuyvgdWMRDj/hhs09yfnB5DjI1B0rz/OaW0
pEFxspVs/2WNSOli2SZWtOp2GbBeZPt0FDlEXarxInZqJVbCdp0/+sHr6BIp0O98nz5oN7qhL+ZU
+QoiU/VSdGK/1x55wn5ODp14gXajyjEjDczkzY37ti07aImqszGKPDdGlAEsNFA6Q7OMObq0+Sei
/jQy3JH/pR7yeaV+Du5v+1ZS429e+YrmltvYj6X75dSAmyIHpsoir1X5diPYJggjBjOCc1uHvjuL
Wyg2W091mznJHAp4zc+yzh+QSy9S2owI0NWIkwDYhxGUjZvO81Y3moRiKDRSEDGCCPrU+hzVQpST
XR/wd2YInworHPh25H8Gnv9i+UdtGV0WXzkB36FPL+NL4oq+dLr/GO+OgxzT94wppe1TYYsfHbkZ
7KKh1zSQtizPBez9BMt9yWa3TpTqz+h+ZQlTW2r/VZBJw2U7OfGOnB6ec7+uQKUWvZuidA97T3cW
NQL+41F97/F4bj0pnIKh4ktEvAgTtzJR6nNtGsqlUgTa4QdSogf1QvlBJvhxpTxmMNM0KMy6WNoS
QO1tJrIR5TV8L3jA0iuPRbZPSONS9CJu3dqreATdXGcXsKkTTRxlsVmw5UA25psJhHMM+U6EM24v
rdv1EDb440Gbl06A03AnUeYUQ39YTI0TohMt2h4CkPQC8ySkMMsrOq6QTj8fNpc1RtI2eByEiKr4
/6vbFp3PI0AA13eeiY7/qtrhyt/suSMHH+UI4gQiWzIYd+sEYIpSH4nbjZwikXxt5oKRrY7SDiwz
ZKrRr6AbKvF3MAUxhi1V42E1ioPwbDJe9TCrMrCgsmnn2wDAGx3xT7DuNwn8+FJB3q34pDyIG3Tx
NRLNutYHAKnW3Q1g35Ss/3wBjqddatZuo+xbXN6ar2/o/wOYpS7l12CsXHImS2uYZOIyDRx01u8/
q91mKDJSR0fo4M7C6G1sHE4hfK1vaKImU22v2jNC8tamICOhacylvYpT1qgI9o3HEymJ+G4L89uC
K0ZcFoAaTIct0jRHPU11dBPE2u+Y4Fl1pHzcc0K2rIpxy62taCv9xiRoaRGG/WihxWOmhzNDvtKE
N3BnF/G1aRfRWWBIOpva1NLLnpORWI5TdRMB+PtYsmRE5Ge3yDO1ExG+lPgLqFKY7r1TndBrGfDX
lemEESAhzDIZXed/wrSeT9rAWQrXq1qCn9dYOnikEE9mV6nLYpxss8MbSoKSD119VsRbM266IYSn
L88Mm5O78wYh4OMxAUuyCe6+3XIu6vWvT+A6pK863XNz+141/h0TDiqg+PuuJ738gNR0aKteQfOS
PqjHQYXw5idm6z/AEYM+0XV0ydB89FaUjThCvttkqq+f7ZtEzACN0Eww4yGjnERbhp5ThgiDBTj1
cXtu72Vghn2ueoQ4Cshl0ly46S+iJlxtnNsgZ3JmpJdVrOGfWhy8fa2pM35fHHUU9m3+OW4pKvb3
Bskdz7pd90DYWpnSTvmifUuwbaH/mkI/dzwCzd5eienARwaWunoOCM1v4gEPpkyJSPEpwiOhOlMR
sTAhGxvwjE2cxss6sKy2NYsUx0lxNJ+bCJh1csh3Z5hUugUQtfQ89XkAkxNrAryv2faXdgQRGOp4
aSCpGmPj2iHv4TyibPd9neMZDXo7s05d3MhBQZb36bV66Uie+dbqo8bnPmabMtqgYquo9i8OYEWs
bBA/8HxE/Sfs7RAgRrGIlOdaUpRtwuIIVpmv2TsaB484DDnFvk4G8D+AaNs/wsGluEWTEvu1NooN
m2heUJJK/CEpQMoXho8GdTW2XsRgxV1hAFhTB0dK3XFssN60sCGP9zO2eLX+0iKy0gkwXWiCo94L
6zpcbsDbqRCUq2/u1trzsMuFkkGVJHfAc8DwGhe+kG/2enuInKIyxX4LSwbGQOdP2YMUxzbKOFrI
930dR44XcBJyFY0bc4Xe/kyQCdaO8g8pBMap+laV8XAsNX9eLGx8QK91/8jFqnuW0pBU0FOH7SMh
fZJ0Us5T7+rJn73t/bh6SY3PHOJV43zTTBZcRnmyzNklcmR+qprx/90p1aYsvULW2K3sDSBT39AV
wpbPP/jMebHFP/SrbjXQivj0qprrfrhNHPq1oQjw41KyZwcnu/XogO7RutF7A8jr3vRE2gnSWRTA
J/9EHKPZUx9y4Hzui78QH02UWHuElpR9IJXa4DXfw7E0rEkXan222B9fTf4/U707NBdYbCluQsd+
R5PHLmZ2NJJHT1D02yUHOPxFf66m1N3F0ERwot93bGfwGGYbVRyEznwTP/J1wIE8EygzkL7cLM0g
cgb//hRy+k3CmCOtaLcrYKmC50rlzB+ZPODTILGgbOjUuEJtHFamLYptjkRIWgRxJJd2vlRh0O2Q
A36AuvHHevc6+MXjOKD//VW+EB4mY9L/+DpR9/bSSQ2Wwj18SwLDfERldhn4pCPcDQVic5wl4pRJ
yjBg7aCIFBEWPyJ38aYDNuSTOIRE1nmIGDiiL9c0GQpF+eLENqch222XUN3L02psKHinx9bY/Tvi
WQUswSrmr5xX4o2ENGgTQFa8mOi5BiwPfNudCilYk6CyDKfFORwWqdmibAxQWPKgiHIXneeTOADx
+B9aYowYQuHif9KiSHeJhP+xvZFJPpJORN8oS6SIIVZpKZDOJESbHGvHJWLah9M3DCv5rcCLK7yu
qvVsT25z2wgnn6E/SdJoYOsFuLck3yK6waN3jW4u4V6JTTb2RHoElEOfJew9YKSYsUH5+3Y3gofS
QNeo/3vBMvvBH2STX5kw0vE3XfLj6voj0t7OzTijZjgdnfX1iCEIA8d4OevF/GDdQ+HM34uewZZq
YOgHNREj4CU1Oforw5+B258ZLjYUj2nQQWt+KalUltFGXBkoxlGSCfoTed87+1FTFpCG3kH/iGMw
RsiKSaZI3iwF2izIAQI4XuvYesY8e0BOOomnzQ1p7KyJ7AAvsGERNdSaosneZncwdpLAgTs4a9FL
Hv786oq75fuRz1G4pMYOmvqn+zauPlkiXiwYq+SRzjy70AZsQcDToTHfbM/Mok1O2fQzpDtMmLKN
wv6w9guvNbfqILV+wob8u+2hl+uqQmAV4MZ6U+FTEFGOyae6QaKVEph7KehKMaDZwx+FvoWnS/Cl
geCMnvtGipUvS2bZURVONVH7xhbCMMsGtTcbFJt6cBZVhvVwYmYaO/hTQTMmWKyeA4lFhlVnlaUS
u30b5kPSKdIzbPpubduOfBAd4PgxmIpF7Yctoo5VTGq2BvXC6D39Iuj7ibJlgbDo0qWVXXdK641/
KJm/0GhXh+O8H+d+759JM/qH+xXw6BknStIMozGNGeFckWwePQYHsfNLcvHsSFGbva6rnFIJTmv3
zM9xNb3ZI7fhMpVTp0sgkVCSSM7CTyCa5EpklbjuU22uy2pF1OgvYSJijySudh58ZYXsOKBdko7d
9n1N/eodWx4kLD6ZQqAvDYNxZ6uU+QpBTPVgncpHPNEYGWHv/HESjCk0MlycmpK9ifzowFG9RSh0
DmgpsuQtVhHIr97jB6o77TBKSg/AWBsPNVmSYxRPl5JQE+B64UJ/RSjCv7CfO6Bq5CxgyQfULOhw
nL4h009FvVaftxK01ufhGkbQW7K0JmOlkleVX+oPenywodjhowXJVsyIj7R5uPv91VFAAcG/webF
wSl9mfTcHF1jlyJ2JCjPP6DtmGvgE6UbW70O6NwoJTvZIMY7223YiDgtGgewUwoitxtuacGbQiis
y0YpAsESMJ+fdnYywYoNvAaA8drBGLq31kybggrmw5Wn4aV/SWB8lCiYQXxjkKjqyimBHA8wQxMK
cRopD2AXWSxaIuhIIlk/Iomxjn4Nx4Q6M1UrPmp+BLAOiZEymXILaqYZcVhLseh1hWgIB10H3xda
9cKQzZ+F3mBee5AI5YIqVqGptLXfuAETjCcWe7A2ewWAqFmS87JemPOJrF+sxL4MvFfkDqvKYhFn
tcvGtMsawznHlTO6VFx5Lu8IWY1Udon7pQKvM5IkqPW52kO7OZ/O8xFBmHif3luiwxpsx7u85EUv
jxGYa5OcEcOKB3+G9sVd4CruQsNKBWR9LUdj+1cabZYcn0r87mCpPlrTNKpIvuoMVUIDIZVSLox6
8U1D/Cgy3bbYjaQVuoWfS6kMPISsOXtlCaLoqYh5K9TA22+co0vj7muG9rnigehjBswD1JgDeYlh
OWxO6mxbLrQJ8z0wNBqWXGEi+H2jMfSGfYTlVMuhN/bT5r/eovNti7MJo1RDQ9a52El2xxpXW+OB
qPhHQjNUJjMNbj8ffTtAioTRwkGCQXxd5NPSm4xdaxoHAN60H+il/rTNjs+NrJhuD3V39w1rPI6y
wSyyyIp5Qf1LalzqNcZPeE+G/OE5lktFpVsP83YrQThxNiPMOmGZ0Gf/VNW7H9WyYK0hf+vwI3FZ
N3z+/hs9/kPYmOaDd3sGt1DpB6Igima3zxAUpevd2QZ4WC9XipX3/bU6p4u7byxCyg20i8H44sw4
Ro1bayxHxAlQ3l0jQQMaQkXEeLENCmPrcRUGGI8qpmSemWsOxcRqovloJ3G7E+zVDYZnLDF1geGV
szlmFCTNeKub29yPeEXY5R4Msibywcyn1Cdrm/hdGM4RbqHi2iITnEVJOk/SYEv0cvwU4EfBS6Gx
gJjCRKavXyhCs59yCZll4yV2koFjID5TtHJZq2aTzPRfMGsoE38YZq+inl5gYZld572VEdWUu7Fk
rOZkuS/1whTUVWnsccTf8AkDQHXQKqbT0fUSthf4ng==
`pragma protect end_protected

