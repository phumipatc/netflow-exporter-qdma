`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
1UDPTdgNitOwVEhKKt8rsv20/PKZK9Iz+RE03DAn7QRwPiqmLonNkIMAnLSjlTyYegQzVhjp4YCz
u1+QWoiZ5fgHW8f6nFU+g6yiWM5tj2iL/Cr4J2fYYUknTdO+cGlbVeAAod0KfQ5KZb8dJ/dEFGBK
6gpZyTWg8XX3cmT57JNLgThRE4YuYnxSZsvVOgZBJgEMsp7ETFkTBwyYD0gcLRXBJ8HCwrIBesdp
qc9W1opVJpnYRif0LrUy5pgiZqWXRbnPZmFeTWZYJDCqJXhIphOQxBUx9QjYnT72lgPbrRHDTp3c
pyXke/w5rtkACjTr1L7i8rg12gHYh2CHtOFYuA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
bNdtXC+LROY5xClz0ZpFlD5bGE8fssYRakKM8wcgmqE9GOvgBmq9O6zS2QdfxXRnJ38XQBQwm+z5
TtH709kKW0CGMjEibTXwJ6bXLEJy2XYsHcOR7UuH3WLhK8E5X4/+NojXuF7EI/pUic1iAMxqcW9u
WPyyMRRas5qaiZOFtNPQogcAHey8ea7dHNHYPY4d9q7905dpt854UmANwGhf2p4gUdF+8YYhFmrx
QeUt/J1oXNz8xX1CIB9sx7cSRi5tgD0j2YCYom2ZH315RZz72g9BbMOTX6R40b1uUNh0YHiKHQoS
HjVGIpiRiVwqHgytjzQx4uaJ/7S7nZfzWlebOAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Vzw2IHQjZlHVqdq/CS6DpYQtBVH1geu2WTNc3Z5m414FXmX2cezJL78+USnGKFQNoqjPlhdtdLNF
6lbpPlNQBA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MHy0g03LLcUo/Z5z9APIDzzbn2eeG7zAHfnAE+dIFavlrAL92Ep9Ud8h7LnRmOKw8Bu0Q3xKiWBj
Z12kidwxiW8ipLvu4u+iT8E9SpjL63WdnzPs6OaOv7pM3VoLV/LFWfkBiOF+U0FOYUbblEHbMnos
5ZA/rOibXtQbeSgyaD8QdvswPLdlqNGEkIeEiY/5sA7fT+phYgIb6aZUOIeQGWI/Vchr2+TzK+G2
ZGs7Ni1kGNc2AM4cUkTB4yUB33S90y/YT/vMXUhPLqzel+ToK8OFEFlGQo6qiYLXuOwmqP9w4aoo
E5fUEQSLK5zCVBedx5moTeBJ2jJVXHZ7Q89ZoQ==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KlxEw4nXQtLiCEL70btJDa5qQGG86PJeFa/qoHRl5Uk0p6NbX8U+K61MQ+95En3cO8Ujrcp+Kzh5
kwCB3waYp2Q2TeXtdRwhT9e89vxiTLKMyx9D5j22yE7XrgFuSy/VMoQln2z1j5YtdwvQv5qULfSk
04Oyrx5chvIqQewVJON98tNLVy8XDoTOKSAaELx9Jl1TdziIVOr56R7iG7i/c/mC/hJpIbvQ1hJs
A44MYg96fNl+3vFj5VtgS80c3Na2/tgnlQkrnFS5DsYIUnpCRu/jM39IHS6y1YJsc84YM6r1dwPV
DqWQnCLcW7iZjso6czJI9bgkYwVn9lFB1MUUIg==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
qs/wZjOIxalg6eeXSLyj+CO31uvkLpdrGhcmMOStrjMUncAkA1j5zrGzrUq0TWxKyI075JyZufoZ
+M+gYdThiBTEdy/e6bvwZIdMvOBFR9VV49jQxutl77QV51WaLo3+D9A6sE8iM8AydxhnrlO+outf
jFlSWgT8wnVVsOGD5MA=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NPSrvH/NwcSIxgs8eqaOIHXTKw8fxDytYnvNZJgaU5dlFv61/mNXt39QSPSKlAS0XFItRNSOhzEd
VTkj71abe2kk59uHrEdLFKd8UPC5vZieGkWIjzBLF5ykyWlfi5cYQb9h78/SjsN83uc1lzddRjIM
+yIVV/XyjwEdLDCjvVnwQlpKXEO/zeCJ86efqD1tkHW/FgAv85msut3XOgMPHOIz1Ryfoglpnm+u
/Gj5VVy52DDF4xgOXWH3TZySmxWu5OpqU1a669vydIzr4z470zxLVbnWeLN0mSxtkmpr8fLR6+Lz
Q+csES5DQdprF/7n6VDuWKQnPPIk1uwen/lygg==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lMs54kRMGMX7lpbfI7DA0tPm+tbdTEJ2sCqER4O+BpwsvdFTs9T5O6kbFX9Qg9SlXmi2WkObvfZt
EyWYaFn7dPGTZFWMdL529WJSfkPeU2fxd5vgd2YVR0JgfCHEBHPmSAsAVctNQYm36B9uti167gHf
T1dwUNEUUbaN5waWDrnCmRjER8pmKBa/EDIVHZG4P+o7gkoV3N+/TLAgd08C+nZ5v8zTCNsQRYx5
mdPbfhRwP2sHtfeK0UVowF2F05WaH4RnED20CV88F7laT4MhcnqWZRjuzJUQy5I4hXqwzZHqWmRw
AoG/O943u0B0+vMN438BXHiLdBJmC+Nx3HlD/A==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
epxDSmcV+3SCPQvEKHoxn3Ae6crH3e9EhTvNZc1O93cT58Yqn5Yt3USdpQG4K74Mk5QrYxq2FuAK
bzmY0apEx7iCuWdsK5D/PWcA05KQrgDf4x+7A0MXBpE8Knm4X9FtSDuMLcKcu/akv5g5cGBzb8Ca
2/0rAFcQSzeE80T/Z64=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Noir+t+a0Q36c9OUR/mVjy+Z+K/86ysgSD1sRw2TsOY8Q/uH1YEbsn7UTd5YGqQrGf8DmMJGE1XJ
lWKK6iZll+zfOY27ywmw3LvGNDSmMd7Pt5AuhglEbA09oG7goZHKeZTDZMLUh9ssTNNKAFOUC+d4
CU3RG1+0B3cMECT54Rg5+Ke7pXK/PRS7z4UwVpmBmlEYOUZ+QyxOdwLmxFFFDRbIx/Hh4qhh7/lE
gXkFQkG4K16j9BEPsRPXBhRsHwrpf+jZrPpPzVW3HbwqLk9D6uzlk5bD3lKChM1RvrD4dryg1CSg
esBlYyo/wy9qXVxjWDATVSVfYftN4w6oOe8p+g==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15584)
`pragma protect data_block
Fr7yKMBKqdICaBQstWw7Z4v9Ra3LD5IvFiljj2KR093AVN185oVZAXBG8dKpMGdQR3mRWGfMA0CP
kDkwJMGJ2SO98yGvBAnygq5r9YH+EvdsbSwjX0PjDtqV9x85GXQQR/TmHqlz5thNp03C23AqCf9V
OoQAk471Mv0SKBnTQfWwpbJZz90hPcVJUZqytNTE4Kk5ByjCRC6fdCdT36xSZ1dueIJEbGW6Hsvt
9k7wTWa8DbmVOXnKy8CynyHZRxwNd0wj+nyywUaeKN27+X3Cfa14vZCW4aX8F1CqMs+FNatRI01r
irZGGkFCoFS/4AQo57WvHDM8hknraCeONman4rbcE8F3LtUO8ELjZHeLvskO0dex2d9KnUdsXewN
/K7hAENr3iozhnzfEX8FwTABrmty5FRkiMO/o0eCC2sxbIjpMOn0qQs7X3AYaiimSun4GDQaX7cN
XLIngnwNtlrX18uWXtT26boMSIk6NSTAUQC+gxdQ+pOFg4JVVIKfk3aujOxsnZN0PeFLQmEOp8N1
OtOUim8tH/yI8O+99sMggbbcaDOFn9TTpzGbYT1tfeDxoOx+nPVTVkkIBiyIe4TqgkHm7vHY0lNt
98ffYOeZ1+F/GYGOcA/unihu47HlH0q5C3vLf+miaPsHq4+qY3o9Iq5B7CApk3KWz8aiu41mJ+ye
wyftI+Qey0MXTA3yOwU7urtOPHE6+CxlGkuR7+POD9FvSvBAdrR/xOniHNumie8BhM3ScVDNSU8p
w/txQ51v9uMLsgcDbsyPJpHNl5qwi+05JFDEpCjrD+mRCI34IMIDbVpS8A5oayTFYF5OWKbLvZ3p
pHeOea3fMKFB19lZHq9q7uEMfL2rcasj8Npdg0SosGpiHUutvMCUc1vOg1ar6xhE78Wij5loCqa0
uruRJC/Hyl9z7K3AEQPvovxipOihk+TxMnsS8TcING2Vf7I0SdA6X8eZ883hwj4m5SOuunUnyBwi
NrLMTuZO1B1U5Dckdm3mabTXFHaf7jafG1L5Qc5qX///t7JqtIJOKR7wBVYLpyvIOT6RgvnAMeok
6p+zBeJcKnl+0SX3BuFWRiimlAoa5RbjTn9V4mq9yjfn7p9S6LfiIlR4nEyphNxqGuHrAnkyExKj
m0S7+QHmW1w7YbZc88XP+LKe5iIvip4F6i5yE7+wQLeN++xokOCQlom/mZL4ohvVKLA0nwZ42EnB
DxhJSIZAH+LpCAnWxfLf7qquYE3LXBjKFqxdtGFIKTpW928EcMahh3ZrB95ZyDjuLpaBXIp/cXQu
6bC1DLt+aYuLXMBKsobKpXdBnI3lBd0mHBbLzQ6Y41IfSFjdkz5W+7TUVxrzsl2Vs5umpNeznzcx
TN8xyCDLf3/VwYrmVTMP0sU8u2jkMhRV6Xt0yePzccL1IC485NZ+a/Mv0sPDQI8vw5wi4JJ4HAEd
ShWFs98MZv0812INmoBNfuxFEjzaOsLa+9Mr1noss6IHXZjwCUDLU/o88GUqDAucTifvxnd96Qm8
aMHk393yXw4l4iy8Ra/PXbqPbHusyvIrHfL1fnTvSvR6ozRj86Y+cptUihl1eIK7MY8IfD91OvP+
7A6b+SFvaIy20pIK9b3GGIFPMBIz0umfeWi9rh7mE6p4/JytKCPyWww+8Lz7//GSxqJRUfLrn2Se
pHRNFLx1TOAEBsF6iKVuN88iQO1/aVG5b2vIOCG9Bb0uhZOHMT9YN2dybVgJvg5mOSo5S6gNljTX
2PkdIwpVw6WfpgISDwUYrSWJNANKW6J5LKfMeNjWlrvvEUD9qgwdtwDi5jQKJ15VXx12AAKkvUQD
VMEEjXz1zzRUxIqi6QzcR9+0R7gGFZBgPvE5JynZnbsxHe8EJaGx5ABls/kFf+uVlJOKYpxI6oVj
ngVG5hikjiKRKLyCEX4KfYTdnnU4Bt9gV0M+fsmycos6s2HKPC0wusQbCClDRqNAcUwomqi0x60i
bhc9SLy+k0uTmJ5KrEgpQ+dQXd36zwM0uIewGjnWj9uFgDfRzngqYbWKZZHqpimTzWEG5SospB0u
xhk+OD/w1GVMJu1KMcFAPhhji5iN5lLSHOOkBox5tXdlXtocISrkMufrsnYBXVJRjbmyw0uyDEht
f8LVnJgT7rw7rgjQfDjXoNbt79CT6NvD6cVI5bWshbqMwEWNVS6E96CKYpeijwSfRCGroortaaEa
/4HKjjqO3OOuVSiA/5IROV/9siUlk9qHrIoiU8mwbOs2+i1OtFJdbHtj3u2u/clmNYBZziEsgIjJ
zb0q5yQuK5SHa/pdfz6L6ZHQ2G6TvBkmwTdb4hIx8vEBmNjCEPQikWJw7Lh4vEQ4osxv8Or/jRAg
XQFv98bkJdKy5DnYT6GAjn6cooViMzDbab1vecnSGATpubILPqUTmZJCt8ERmUvaoFE3UqRvuCFX
G2clZTyCDfObV0B2Htogx2RyqPPYiH4ifGNJMTcCPdKDlloTpsPvUOOGQkFCPJcQx6DiH6hHi04z
qiDIoakt4BZXsrfRoc6A7d3kUL2GPpJYAdnZz/EpOYcE8usM5XKCvk8auSHrJyi33U3vRwHtyPqd
tiwTpmEdj/fbCVk9nN1G3zUd174zjLp8BwHxO9Jd7TqZXjt0uOZksG/ii5XWA9e8PSyHeN84jRFJ
eM+zKnGWpzNXSPXVU3bTB5C6/9srNqk4n9aOUj/Amkr4hFjO4PAirGE11hLFnuDFlK5Sn0FOdvIQ
K96MtnbYsU8fVura/l5nqY/zB6mQABynfOJY2MCBVRYdl+tDlviYOnrr3g1G5UqOhrUSsAuqbzc0
Ift20OrHt+NfUIbUj6QEA7D87FvbTUbvFk9zcSqzeuEFYVZVByklkdbBx3Wy3F25y8zlIEa6sFmy
hX+QlxlUMaULabmMRHEMFBv1LGJsQ3M4VhAq497ETyDTrLmaiE2PLqrHg2EZDi5BtWsf3p6aBcMp
FB3rJesq57Pc0w6tV0otWXxDuWj3mTRao7sr8MsHr9jlmHOaYS9NAORm4qcO0FJc50HqEDsa8M/9
7kZDIHhbxCzgelDq+Jci+Je+pO5jwCXy/M11DF5/gUUgYmCqE3U5VpGJS+ir5brPxUEe9eXYBtaA
jr5Cvo76aKmt2DPRfBBvHrEDXlu2Rzz0i31dD4WkI/DDvyqLpeOE9IvkFcp5amDn/Z9gOzQyX4IP
5qSHRO/YBNsUlBtBTHODbcmKYBk9YJ6P5nyOFwKyPvjlkPmoKbvBzNr17PgJCiBsS3FGcc3hfGfA
OfY3M0/8T4xSWsHf9xGhmc6v3DbTpC4rqLb2uuTvKRc4msaQmPGW92PYb4+9BJZtXisiFL/8gnXs
qlccw5E4ox345zPiSGTo21TaJTb7fyOMCe9aS4b8qGggjjXsF6lzD1yhUk4A1yYcPO2C3Mg1CmGz
J+00jnDWFdZxIXx5UjkxNGddDDdn6qnL3a81Qqa169lmkxcT/kpHuPOkQleACimrgm35ZY3FyWma
XXMy2z5GsXtHr2sxKZrdLseHOZFOCbLtDBEpwBT5THMg4FxrDoMkBfqXbfBWpE9ZW9+diEXSoT2E
c7dpZtvcqo4kn+R+Npv5OgLWmO3N5xbq6NlfA1qHB2ZL7gRFtmKi1EvdOVCn/zQeWowu8X8mYVPq
GcSi4WYcOqbnkrO5oWc1BuRNlMfD+7oLhHVsIMSJ+LX+WV3YIiJdsThwld5KI+JID6wi/57jq0W0
HCzjvc/9eDu5Re0pZJMkOxzIZhINWjzGJLk3qLENIqVS+WSiCGfbg5zhj5ngdgjFhMsIVUjubXTR
pYaH/Xl42mlxd5J31pstXhspZ3363VUIEDpq9oyr5ML2TIiVxsN9LNayMmyUwi7AJoeRQxqZq//a
/KnJ7eR7TPItzssZa6G9MY1X2xA+FUsWJ07BeBJOkc2M7jsIydggJLt0a1SpCjIZtyfs/aQJehZ6
aD6bCPujE8VsgVGcBblECi4c574/ss/HsUHGzVB6GF3O9qhXfHGKDrNZBZxCg19itwatUf2iUoru
sGpnzLXNEEcnzRSZ8Jn/21o2a7LMGxmUG+CaY+rIGqw8RMV3FEc8D5oN/kgbOcaSbQrYgKxGUcD0
G5HrVZY7359faZHxI0v6vBjXTzOz09s/CYkuBpP8R/S/usdQ3/pNiND5zKjYqU3mNBRTuMhl2ule
7ERKDLS2lPnjfzi6yeRXkFU71MPeY4hq5zg1PkjhEPUAh8F7EZUq+2FUnn1UV9c9CRQrWhGbvfKr
XaXkColVHUMFwej0hTIUD5VRmIWx2zwuzb39AhxOtUYnPENUGR4z3ZHachtzvrEYLSeCP62wGN6s
FcGiv0FJYc8DcMRkAezzrKfzPS6kuWZENbg7KIHnrdoVJYfcuVbTKM5LcuCU71ba8ro2l6I08dyg
q1Z2GuK4H//V4GgsR5+lu2Mr3jf9b/sVDsRok0eVNOuJcpX+gyE9lEa6hZJyuGo8xme/gedf9ZJB
6LMyNXvTbS3cMvM3t7DvVQEXs5cRYiqnKwtceENV2cKklAMI7kMEVE5m8NwAR9/DsXBpqxKSe7UH
k48o2bKlNd0QvgB86VhNVJ6bufbL+m9ovgJj9G85vDWvSDkJ/UCrM2Vb/UW7RnSrpN6l7BqarirY
EA3EgBobMTmdaiX6thTJqhqvwZaprLLVOqaPXbPOQl0W14+9eXmAa1o2JlS6QvRoiB62Vnw0F3E2
E+IBzFPrdY4q6bJWsuoZg9ycnul7VUe+dSRBQ/tSj9mD6/2zO5V4Yefu/ChdVhPSuRz/1JVj1wwp
X/GD9/plhmcGku6fuH7C05GtQ9a8dnkVj+KSHLLOndSNn+1I4lN1yVQXLWisLn71p4u8c2iefuv9
dizhxUfpJh+m/NV+dGYm9N9wpvL43iKsLxVQ97G7dfVHnikBKNb/kjwQpcaUJgVveigpASZoZDU5
T0+L61iorLHUBC5+z435XdLO6FHorDs1zF/TY8IdSP6EEHbNuVrWiRIBK1g1uuBwrNcMKCJJSiqM
1Dp7YUGc+3RClE6LqLQZ3Ypoa4ic58Lh4blmQyDIzOkoHgVYEsXIotjujuLf8QX9jDDMSxZ4zg0F
1qVL8MBRsmRWibXVj+mJePLrG5sWud858sMclFS2v910Bq3ybkuZIY1vy7zKp5CuKwe5RZGRQJnU
WgVwRUgdygwK92HV1gTVrmWAID5d+qFiyF8f1L61RqDJIwkCgyhSdt+vC5o7cAbqfp+hm44yXxgG
IsHKfuMIho20cilh4jhr1j6y2towcPlDzAhDBjVruKigg6gCDy98keY0a+ReNCUNV2gkBEa3cxZN
hQbe3H6bw46NJ3/et0V4LAmzD9u8bUtvtjBfoV/ciH1CV3EVkfAIcuMEMFiva+u+dhksMoXADRVh
bOYNAYeIfongYhe5uHLtxlxg36jVAYpiEe0PVuKhiU8odSb8NR3gKF4M9xWOpTpumqsl3bQzgc0M
7rrtjLQEi+c8+FlyaDH8ZXm/sq2CwFBtbk6iqwPG87ENujR1VaXTqrokns+/m5dOmEWxK0l7O1VG
6XGZw7mVGzIsXDfpgLVcEEuGIE9oZUo130Oz63kBVQ48hlTCmg8kVxZu86Evcdw1rlE8RVB//D4g
5BmwrFh6tL5+9OhUDu8iYb7EZQ+JdNlf24+hSdeeh7xbGkd4kL4B3cSmKy3osHst6Vl8ExRctlg3
ie+8i5bsQE2gj234R2A6kUtd9pYj5Y8vSzXIcBEhpKQ72j8owcILwCOi7mOhTWFCNs4hhMFfl8PG
LjfCAkGG1n345vNkFgj/r7p3/uK6QXONDSFzd0Q5jCJVz2RiQxzm0NUqVScG01eQDubajRfd7BfY
af+Uoiq6JCQ80TSmeIbLYcpBx2JJyGaqnh2huuoIZLxkYN5FLvLk4qwYO2JdZlP8OAgjHhT+njKm
2lQuF7MwR7EDC8aip8Q8fj0TcxqxvEkoBrsF3L85d0KlPs0YinS52K0lpYe5s+xtDeIgZk/Ibii+
FJ1fYJaGc82SCDPQE5F+OHabddIc0hIvup+IDLuqRFEh+NNmwljhQUT3K+pwa453qDndQI3EKtNA
IzZKHPwOprxvfOsotb0D/WrEOwAe3pnzr1YmFf4f9xkh9NflQZa8BZE4/1iZ0+/tX8zm9BH9U3YG
6g2Kv9seUkhM85WsxPIHFrKemezFC5UGay+a9ZzGoC/CU8UWUTHpygi+Gx/WaeNw/LH4eKxGrR7f
hbqzYkeVKwa2EvUYRewapzo0JGKeBIBd/MKjhFVC9doyNEZwhzFyv7HID2OApJw9OaJrG8fvf0Zb
INFdvUgImVcIT3JaARwOJy3n5mKehd5athm65OrwW5Yj6LuYJK0I74sEi6gPkzk4mi9z0jZytH4s
0NvCyvRpOzPwXQ5UVJOM9igZwnpMNV7sEJazcf/3/mVnGJVFhDssYJXmguUHxC+ngUZmJyevp4An
GoGg1HQqtqCc9DbZcKx26EbqVb8HdXtvpM/9x43cxfYUkTmFLwq7k2IGstsf087hx2t44U59JqiE
8221VNY2xWYPeowadK9mbGUuDbZG2EZJzKf0g5RScgZCxYIrmLJfaMj6f/j0KJ/n8paPFU7J98aN
Zr+b3L3wZaYrYWtg0p2uk16tZg+01mxa3UDXL7WFckl+lti7Btr+1DLPbAE+c0k3ut/l5BTFmJgM
rjEPNoMOk6Us4aD9teAL3n083+UMIh7Gc35d+27kHbkihx/Djb8OC1CmWSVMCe1SsVcjbjRs5zVX
JTGxQsS/Q7ydhJJrLPIKddhnjiVwLqn/WT222fl8dW6XtmM0zFga2nCCVAkR6aAeZo7AqI8pd4bG
EH2eaOr8qNFExI6fPV28ULaY7zQmVO2JCa9X5lcPzVVSWzecvfm12kXNp2AHtxUbstgZlh9AwGfA
O0DiHzUUs+I3N5quWp4zzqaju5mF/BuB1KOsq5qLeiz5QCtDCpwBuMdQ5fLEoubN7qal2QMEPj3d
n9vKYYLucfmBa7Ba5W+y0OkhvgNV7+ZzP3STdplNGscRKXcvjbS+UbnmZW/Tu3JVjKgqJdrlikXe
R3iSQ81eycXRIc6dvHTzrq05qnveT+JHC+UQCe8w9kDOPGSB98BkbRDyUKkRcQWpWJCMDY/wERar
qBlOq9xvYWmTVtccKR/DbBeU0mhsYpTwUAEzhEl8K0UcCT7p9eOR4pMaTQzQjRJlybqulMTE9bg6
toXY8OsOrsJsom2tLEOogcuLAx0Xv5d1jAddCVQZethCCp7XylDMka9XUWYB0XR3G3CtOzxbd6Du
DrU19hlpNs+gwGZ4rqL95/QWQRuUMeXMFSc6tV/fLtPYx/JpyM8ag38kjWCuBfVyRnrLtQtRmNwk
pPYtG5VG8bwAh6Kfd/LWJ3/ZX0SqQzwph8ohNLMov3ENCdg9M3cZpEBmX5jDT2kbXXTqeu1zJnkS
W5dbzIL3ZA/Eulfyg8IJ7UvXlSTw5tDAbFoFHk+G57YDQcK3CNH/VP8psel3CtOviF3YOz/A10Rx
0XeKh7CnM8L0S2JcRYg+MoJ4ogz/s0JZyaQ57XvwA01u1J4YJK1LU6UJfqT+ooS1FpGvWM2AI/2r
pLMyFOgmk91HFMFAkJxVjEZAn2Yin1n+2UsKpEd3t53omBdEy5OwR8UOoYfTsAcmHuANe+vKyep2
Uf69OavXylP9e7DT32u63xhOp+jgH9/lDTeP3t5iuPQp5NekHWwniHXedq4O4yF/JqUzd0MNL3RR
nLZzXkUXUmXh3buGK0cv1spgLSg+LUj1+f1UNEPRzBVHX4h+Sdq6Ylj60r0w1Gjy/AGRMFFmHliO
iDBRjy9dAKHeTiI0YQatI6tztwk6+czq8gb1MJxEBEgtCk7q5/gVRe9mq5fhpBS4QxLv5ovE35xL
SlcwK7x1XxZWU4bsS9vN3QhwprVRKa2xILJtOuwQ02O2ddUY23Pq5XIUkhNf25l9ETW3wDNISClw
xvN0bsTqYXlEZs1KDRDLv+7U+I2oCaL0KrqaYK7BxP1m1JlhvsFOXrOO2SIlJ5vW9biOqER9lWzu
HJNMlg47XiUyaIJZWEhcyKtRGq7H4YLWBKwhaLXS3jp5F8lRfJtRfsbPeC1TiGJTLAIO5xb82Oqw
q5FASqzaU381XXcLdW91rAQZbauixafvNAis6PH5EvFP0+7kykUpTHxFe0WJlHxMCMyfFTppCHsf
BwUW2+jnqcNW5CyN8LE12bU3AbwPUNAAnoKHthVnMgv8jNAiVoR387UAn0z9nwhEuq9UfE+TjNKF
fjSDuqurpILoU8rfxbwzmTm4IoYTHSreAnKxjoEbaPxNokWu9Ok5TH+5cXvaMqCuOMcvJhyEQBMR
MYSYfIC5npw1d09ZJpjRfzf0MMzDsXyJnqYUyp9cGnHNx6+sR0iUInyPMeRbqLF3iZFY1rc516oN
VqphDBnq0AL2nRazz6bg599eh8igTnqp8q6zd6EkbtuVPtbc8zaTxTVo/QH6er7I3frEUNjg+ikX
dFkWxpA1J2CzZA4f5NA+mb/68rYo/O0fiEeevBeFAbiHbCIkgxeN+/U+gnNyXpWXmxBstG2lDdkz
Or4XjXJnDyHYMoYexCRhursDG5YPuU59bfgFhUOQgUGjsq/JcxZlN3jagDEItunCOA9BYWSLsjFS
6mqmzrtP3hOjAb4LMiIWdGdb3w9HuaHEb4GvOrCdKgdfDA5n9CQY8xcD3cjXihlsNN1GDeb/i3ti
Dpf6dvwsasiry8LLUhkoHRHXwRpTxhY3/VbLjkIvyHyE/wp9zv1ZWrzYMbAwNOEXzJn/Vyk1Wrig
kpS5/0+36i0Maax6Aa+nrRbV/Wi20DgePaTNd6zaDEVE9MURIZZws9DSVSqreVe9YGTT2ZlQ2t2/
XlOmay+hlaQiWMPKg3dQhscwlURTT4qi9cbOtcnY1V1DhJ44Sxl2Fj8e+55Naro5HKhMmwvHS5S3
/CBXOVjmnwQ8TmL4xP3UDlguk/yEbHhDXELpV93+3U9PxFiMj7VJgxHJzMJFLNfRk2+sSg2RqCHZ
g0p4QHHcp2uFTHobkmkK14U5ZnDGR+r273y1jBv3jLkuXTsTl/phA8/WuTTSGs3Iu1C0ZB38lWfS
N6YhG4UmqauYo7KxdqQ4kGAN7mqcjrGQZDE5oqVUv1dxrboEpKni0rMEE83//cB30RyyAMaCbL5J
UwhRrlilZ006xk8O2PA9icXqd35v+fVxdWw2IA0XYTSFRArdGR1750jikh/dyk19Kd4q1sfp0YgK
JT/Hzu/feIUky6bicewFJiqbe5mK1rOUMDmaYCHo6zZJA5cJxHKN/fLAqcmLGpckmMwEc6aM299I
H2+U4WLhId89mSA04hGVtICzCLLqnCjF622X/SEnf0+0f3HldB0j4AP33e5VR3kfn2P6SqBj8jg4
JrbE/RrLPoJ4mE3AErv4qTeK60z2Y8/USzm/MSb9NsYstL3pBIkAt8rgPEEbUev5KrZOo7O0IBJS
maN/j8Bw/srzDn3dQbYm+X5BhzAXke1eJ7FqekNPaiQINJY43OEV01CJUYSDAMn5ufNZB7LthZIm
XD2ItlUdOKCWlVmDuRCNvnsF/IJWYeqViFFTqdCmFRkIBz5c0dm445glSDcIbZw+I2a5TtkCKqbZ
G9wfLCrqEKfnQV4/OVnhPltN6Ut8l9qjkaT5cwxy49rySbvdimyrV8ft2HuSUa3XBH1DMs/Pez13
YHo8dUis+2mKWnZivs6nfNoLyKVOgEg7G/UVTAhRSYadUBuT1gMuiPo+vzpQKT2wmrpXCz0lKQ6p
O49p1lDU9VwylAL45JgYTx09vtL50kgvPBMNp1DCYeOpPzdd86S1GIYR59SWIeOVW/bBY20NqBTU
jmQJCn2b+voq27oQWLqdLpSPX07IieqEgaeVl9mgl98m/k2XEu4J+ihhmcwsimchYrBGM5iJqEJe
y1nbjJEhHRVq+pljZAAjwOX8/K8AWNk2ofkrJB9pBTrULxJLB5T5vF48h2UOTQWFz0dnbag6Li4h
wPTFrchbPswr9yZr1OJn3/KJbknJ9RV/3mSf0Mh/Zt7cHsYLE3owLa5GZJKYozRpNkBFYpw3BZKR
kz9nicFRJE2/tOY1+/YjjsyASbUQ7omUhz7mobZqF+Q5QI05mPC/QFblsGcdmU4r1iAZV4j/tXNA
67E0zqOHrPsdNafCraNKky3T7UdpNtt7W11p609XrL5D68a0IMhazTuhmSFmsFe42IX6zpq47VB4
M+Rh4rRziO2StfVLpPtg4M+RYKAl67eohfWONDDuxBBiqah345V2YJ31iIJnX05OuYWHwWzeXtqX
UjDYff/Oi1EfCVwMhzjm/J1vFSYwmIknseb249odWOs02xWoKyMuxqSr4h3e97YlQUibE3ziV+3k
Y+nEyrRgCWU10HSCTXr1Hsm/+4pspf0nVhongbJbThsslgKZVS3cvrxOw55Hucfjuj7NYbQGX8eN
lpUVLQQc74aIttEhZho78CA24fk65JoYLvgkblLdTUio3KpMvWcZRk9sm08HnNApblJCGsQ+7S11
16fNRlxt4GrBI6upyCA1HmiyZ70kFG6HbB8BCjiWaZFVEpTbscArnScUdrwsF86VU7cXVMaHis5L
51dJ0rhziQQqVaNoiiOIXmpPrbtPzU0mh74YsiasvBFoUlxOvAUVKl9Tfdu3usQLZZL1Do2FqVOP
h8vQ5QWCdONaCmpB/R9tb0+isYhac6BVUJA/VpHa3V7tI24z8oUiCHdIbnsU18woguCkCNnTGeL+
jwuUqsPP/fGpZDGRlgwn4VArIE+k4BV6IDTG7MyUZeEUMiYjBqLZeLb1oXDRgN81oy2x1Rp9kIfd
RsPrxPtoOZMQA+fUnQDZums7LuHGCNBgHSvZ3A34nEOlebke15m0I0m/sQPJ7y9JCmHxEojMzdQY
g7hmCNhwrASuBOg2SYEnuHCpqrK+QpHSVjkD7AqbdDmuwLanY7CkOXQP91Js605smZdZN+ofrmuB
39A93pjJqR4zl1cpKd9B4CPLU0pqxbZnpb04xUiePLmXnscdjGxzDZA2HW88sFofJlr9Af1LaX7G
XsqEKA0q1HMrp8Zdvvpr6cix5B7X6VfND7BZplwGCFc/mcakZr8H1PSCfQoANPwFCLXVxCAUWwvE
9j02AS00SRWMwHXA7iUuwL6ShkBOehwcixJ/gz4KTSEcQbLTFsldF7OCL/aqO37pQLClA52ZFKHj
v0Yr/7ot/2LdZVwSPye/lZvhedW9Au2f5zcV1xf8w+ODtgfZI/OvM8XKtFN2KrP+PEQ3HEAjYwuo
UcNfFY4VA1RjqNjyX1mFH4TN2bjcrbM4f0+etj4VSLwnOdxITAz/E4vU2vn2Cov3+UGpvLgnQyll
WPK6Mb8F43WojGt8D5E5ZKVNndnxSfwhbOh4IlCWvJqXHnueNntjG8psCSOuq0J4/sb71IGz7YS5
wH9AmWL/z5EN0hYF8ykTXHcYyvA6oG6W/YuZy2MtYhm2v8FSUqXIGmVSzNLiOfzmabbHIzPlqYOz
0us7fijJtaSh+a6m2JCNFIUfQAE8aOzK0fYJX0uTSO7JqX5lNLVpiUQwPgnWJAjT9mWUXcP5Vn5i
mI45nAWQek0A6ZjWKKPVZcXG1kCzey+VYFz2cn+TDhWzXTFT3CYAjp16dI0FD9PccWVEloFX+8i2
m7mAtDe2HxnwZ0L+zBzdvX62T5sgJ22QPRNUfW4R7Z9qCknoSr3fNLETbIniepQVYXlqkkMjaF/U
EToJLHVCI0LSvgA0NLw+ns/NwU+blZClD+0XZmWtecYXNLIOexrYJcy7rm8cRiBCdiwgf51EXpHm
75OL23A5xN5PE2EMiFBMFV5YbwJe8r6p5ZvwBM7WHoE647ar9wIReI0HJyU1qAkEkPxzeEM2kdBK
6hGHGTZ0S1DzbKj27ORHvZgwfCZdsHBsXCcsJvs//91i67QQXBpTpTFC02PYrBJ+497VNX4XFkC1
XlGgi9vDIBK90ZYMp4ZR0mo9TXR1adXUBwsu8cMxNpA+IxI5Cea/trFgOEm36qsSooMBYmg6cmD2
75nTTcJDPE5xeH4rgN3ga6m1g9zJ8kiHWIKclAaaZgk9x2VKqp45DNJf0iB87ch+Ulg7OwxrwGQ4
21ucyXA7QwMm5l8CfQcQiBL3em+Z6HJFSrYgCPpRdDkIvw5QfaPF7ZvQtiSgI98GNnMdDc+PtTMS
UOAljV6vCNGxQ/6PloG0UkFIJBbg0IMldK94yrq3mhZ40zMHgjbWgvlAm+6MTRRCZbbpOB2+Opgk
vNyUKIj50jnPveQvfFpNO9u7afxIkQt4ZhEPTXhS46n8q2gIdLv8ZfjW2XLXI7g1lPYrsf3wsgnh
Ts8Fh/S6M2P/0w856ACi+Xsxx5vpBlumKS4MAM1G9b5UjBXgyfLV9612AoCf+WqY2ZtI0hNxyoJ4
/WM+UaINzITr6kGb5gCMpBIzDh/1gJVZO8Prk7MUkgrx51W8Sy6LBbgSG5cJoDczh0OE6ueDoXTr
WMqrUoKjzrdUznVmkR9OJ1q3d+deuGwmEtGKSrL6XyZISoG5j6KB9WUvExTEIDc3xUEZ19j9kRPV
aUdqS+BG8C217YzXe2g0y7Tu8ObkVg5qtg2wOrSOPoLqtdcsWEc9yGD24tIegixiYujmNcYxb+A7
0v0vfvD//E0B3wZe2WziL5Hilt+5Vy2NiSkouKdR2zNkbzxKfJmofiLGIgYa+aeMRDO8cmWHs4Y4
C+Pnr98K6qy5pANIIEH4s7KJPkAQmOCJ+EzW0ptGXCcy/hiIDnWbocnD3ua1LPwUc0feAIiEhEWZ
htBgkqV4TjptqQx4IZsTolxBcUJOPl6GkAbuZtELkfIMGD/cpKRwzeXETMML2cYrPfHRKMlTIJob
MPbcB12yjKY9NC4ufuwN/XydZiMMZWYUEQwoD4D7eyW9kZjPt9pTEegzNwg8mKk1QjXaAJgz94jI
KWrzAFfdj0EXFMeEifdV345IA2x9awV8KWHfL8ltZDLjlOnl8DfiX+tE/aUI0kZ8wYxiFlxTKTyq
UCSn5V7g5Sj3M85obdmXtCptkSH/rlunQ2OQ9ZUjIUUIV1ekyVlWTdAM/PqBPXj+kv8f2Gm5faTe
DBFvJmE32gkeXfWSzXYQ/ecfKrHyDBT1k+qPmv5XQwKvEHhhWBcWZOMQ+TVDNY6ukdgHn+jtyMyb
g/oLAJwbSNPwu+fcUOgiSQkv0IKDI/n2c1leCdJ7FvggnXes3RC9ESVUBRIMXTfkg5IHiM/WAem7
8eVhUtnZzYNsds7lq0gQLjW+8F6PELu7zGtZ6VLlStGEtPUwC4W1U/3t38O41qkyQmcAgRsnqcoM
2KTIS0wC5i8LfKgEgAPCG8FuwTR7MaCFChHI3dV4S4qwGcy0drsBLoxz1MJKD9mxo1fgkg+wvmXj
3FbyF9tCzzfalr6wgmlq2f85vF9y3v8IdvPg8zCKQPyY+oxGaMZWK/dUhC2daVVaSIxqm/IB7IMf
HDmZfCRT1/GBAqCt/ZTmY7hWMPxEvbkWA4B82FlFmMQzbn8pAnbkgC2L2PTowVWhwty0XgqeVxBT
yV5+a/91P73ygx6Dv4F7AMuiqHOnYRm62XGkAZwqLIi8fde3FqAWuROkVWvMrxOaUKYcCD9+x6Fe
oFoUtU3WlrsJTXKx6wTH53Yy3iYraKrfM4kmD1Uy6UOh59n7sYIrAEyPN5OrUXThQL9lBC7dSK9i
nUpdqAXAIm+Ryjpfu03kaPuvvwe7KCTW0495ovvOku6qrLfP67bbUa7oHrRRgjLReArwk//+qE+I
CPqFw87DYgKkZJ093NBWNgk3JpxetBDkSh4WgHGv+nvCqDnim1X1G0ln73T5acnygMcZIyoLMH2B
NOBxz29XK+fuE2GZoTFNw5E0FmwUvhnJ4F+sdxr9OBXvq140XupQt4a5/KWU28WffpiS7NARe8K8
pT+sIcrnxurKdp/pZ5VD+heDvrwKo1xYvDX/WiACs/bYBt03HUl54S/UMzxWA1huIwZq/PAASU8N
d12cA1IcE8H9JsVW8Bno+Tlc7CQ6E2B+vLhd0mBQqhx0yPss8zstjwgmevvh2fCTzJjzKHWxgxnk
R1DvTjBLbYPn+Vfn8HkM9ecqV3qxbhvfD1MkeSx5XYCrClwEse2Tg1gOB/45shmW4eb5jMDFhhIC
Wy9e9Z3SZVKdwwjDEY/cXIjV+Ei4rfdwqAjJbwI2I1fAD2SIGa1Ygj6dH20BrOkEiIse9B7EZlKE
kQEYVpF821cqU6aJN0D+jEhX0/4/Hw8x7neD2W7NoNTvNs/uCUv2t3R6N+MsH+JfLMu3m6qNEIUB
V/l4pDoypiEDJr4t/I/nI4CzXXFtY5kTFvJl9XqeDqoqKRPK332HhigOyvfJRwyrxbXjeW5IkjdC
S1KOW2gIpaNH3wiLOBPJGNIrk15Xu/sAtNcgy2EtjWJYzgyPWMniPccWVJcQx8966sF/NThgN4hw
NfjTUAiFgrOWUv0QZO+khier6VlSppzJSptf+1dzh38dA5HUJyIJpQmbtu/OMjgTn51RouQ/TmOO
ti/kojypIAmUxiB5U0u+r3EBSyuqlwzRSQyBIq8CCfVvYz+Ya0vy7H224nBHLSaJJL4Hn22VyTWE
QhlxBn2fw6QQ1LS72hLbEkMcQ5P97h94rUMIhkqnAnkjeu4BiBXOnSUZA3kjFQajbcDzd6gcTvXR
eFmynFND7QJeZeFmNd29eCUj/xklSGnbTxsO3z8c1YosRe3HwDKRifz+h6UwRgOu+VRoVbMf3zZF
pj9I+1r8hTI4CX4GB3wXYajLEnu4HS3BCNNUq7mmHsCvk8xIX9PkPesqyjWzjH4BGmHrbRGXUWtu
+6KE0LvHZeol+7yS3A36xCc8uSjGA7bU4worF+645HEZTXY48CVVSD3Qhb9wcn+ZXNG+EY62uXPO
vIt3F1JSN3oyuFc13wi2ukjvyHjc+BEILu4OO8WWgMCxVb+fAdkGEObjcSIiihXJesogEuFcP8NG
Pnfa95QBLe287bv2jKXneMOzFXV1ziyeML9inIMKmnR2tF6utaKAGe+V51YBToqiGEFPrZXfxbAX
oXNEri+ApyNNpOiTrizvAZ1IxjNUp3eClemmgzU9KxDVitBAooOHuVQxdnnACYiHE2SNjEJhxpAW
gTxs+k7w2a+B/thvyiy6D0uxmZtqgMGBqM6wgefthM34ykl9PLUkkrfxNstZoFFEMKwjJcoPpLX0
vHqAcDUTx4yYlBYKC3+UV9XrSijwKT8cJltmrNtnCfMZyIfYyUVpu/Avdbp1YhqDaywZp1UmV9yI
wK88eoTFbVCVyUy7gOmoMG/HOIBPqEiIPYTUUa91SPoB2knQuyCCCKd1f2x7WI8VbFuRjuc9t9ej
3uuj+8RPAev46ubL9l2R3gNngHGV9QqHYMjxlLHDnelW5A1e0UG/J4TgIK5RLpkh2eE0bcVwV8NP
FJcRN2Uyb+obyY+0D63TAxgl68HEHMzBx0ZffyX2yU0djFjsHi4BvzatLjh7JcL14+jpfNzNIvUI
J+5KQk2tVVIgsyuSnvhH/iIlRPXAdt/DVPCGYI3N4O1H8CdhyFWHDPMyBH6YMrzIK3C0KoB2/4ld
ig6m+ckrgNZkDbZc6Qlmsm3nKFSztTlQ3vN088Li2BFiVUM1Ru4jCVpQz4mmaYjcCz2yx7mzFZcs
EuZUqnWOobM+pF5CP6jPjL08oPWorFPoqX5/8QGNXvBchoaO+c4FU0Pm49bjCmVOvn2roEgDdz0d
nNcBMBxJk++ZLK6OtCrT+cmTf8nn843YqGvbdnw53k+RN64GrkIIx7HkN2fAisLCngmCSbMe19dr
0DaotR7a0I1kBF5IdvqaF6JGxR6TKG6LRachsA+Dh/TYhpcpSMZ+NuD087tuHnLLOWX7q0YlsYY8
YsRu6EhNHyxy1VXz/H7h67z7PIKIt2p/pgIk5tgKhChFEkwKgx6ZwUJR3GvqZUO0cyxVV2G7sJTa
v0yzjN+ddtYto6dswu1vCsR+5UPJkkBtEwl57BhFZc4EBj6L2aESMy2TM7QHdIITf11QkZlX+l40
zKmXqSz4ClVg9hQVu4JjIx4zPNcmacWV6vyUJ+aCHyHJ27kSQk/ywRUEinJuZZBWvnUOI1saQkrv
oBc8nsxdiegneEfuX9iE9HaUFvr6rn8WDL9cMyp+WfxbiUTljsjtRVJLw/Vundp2CJ+oeHc7EVIQ
Znyulk8dZUJIX2i02mpeGdPmW1z7e4WZMSVhhKUh/XFrgawaKLUyj0c3Nwt/T5zdu0y5AH8bLect
uSwUWbkO6SUnqxzJB55L0Ko3w2C+0zYDin7ixHIDSCs8vU++RakBMtZ5bGM8Q12Un6jkzr7k7CvU
9CbC/g7q5fmLiHwwdrcPkraxFgylujc00pvRypSTTbB9hRLbuthnOM/DHEQOOSwOanjySA01sNrI
+37Sg+O1nZ+Q2wjm+vbfJiE2DpKfBlKnFyLeKHmMl6TG6RqpRUI0m58hDejkR9CiuyI3JEN3ZLh5
t4dQ0DZ4NT4y020Kd3f0UgM82Ofz7qu8STjnURo+Z4Wx40wYrtVB8s9hOfL78qIAD1AG9uQoNbTX
nPBe1DDqvsOUUTFwOy8KTaFJBnRTEBURoECpQWmPxqmZoTRGtx7LONkVBjNBefN+3wWJ7QuEFPyD
e9QmLotzn3l0VfGIwPkD1gWYNOhpwyCEqHMGmAdYCW0mfo1xA4a0O00WXQQDaFjqJtRtDfGn6Enz
i51mWt2OYtJcCN2cipke75UMKZM3S6syI4DHrsnNboiItm1ZoBUTuxv5kZfPDF3WOzUFTpOWhHBr
8DSfrXuetLRgSyHvr0Yw6g/3HnZxH+DzXzJJvqzt0qDA4m3VNot3Njop61LeEAQUYEnAnNvhzIvy
mxyFoxsWf2jhmuAXdLgQkE8w7Q77AElzLn+ZaP0p5epeJwj2cKkn8UvkqlnjnUsjDKbBPm9ddCU+
3kGF+vW8qMcHaFdd3McJsYeSywGI7IR1mqTQi78Qz+xwPlz0nnO/kTYUWzNJ1XPLT5XAfaqUvyAG
En86nelJq7JcMpUiS/RzgzSdvv3z87W1Gi4cvg6ayRXczjvzBtRkykGXcVSCVDOnxlOTwRl+kobb
3FNT2cL9s/tBjSES2BCE6wFWBLasG9voWJVVEQUrDSNmJHyLRTc3+LByjDMcI41IqvGc6VmRv74W
OjM7ZTMbyEd3GzbEspMs+RWDCml5SZOsASsPzPoOSStAcezgcH98mC1tZtsjSsBon5hA1zYTjvar
AP7GftkpR0oYUc30No66b/vlf3Rt5S4gka97Chk1/kESRrtGDnutn84QOf8khQ97zWUddUr8Fmvr
5BRENNLQguJQXVmKkp9SPvtgOoksA3wd1kJkRIMADhPMoOZk1Uuutq8NrRHww4/te4W+ejwQi7tg
tdVZxm3P7ZpNFlHRNSSOAE2Flq6V6+El1xLXfBBDZk/t/a+RlibfBEy2nvokmo0Ci01Wjo9uXoAf
4t7reCHPYSWtXPiiY11EuNwJDsVmIoHHHFWAK3Xju2/JbU0d+bWHJNvp6ZXidCksnbFACCMVkdpc
pnByaUxgO+07+/1L5A6SvuWHBhEYGcO/Lsd79JBhJ4mi4UCJwsFB6zCZh1gCpB8XdtIlpqdlXpDy
bcsNVPyBiiptoG9n0JdDP/MrvNZVHpB+7phwngW+jHD4ctU8AC/b3fJFu5cR1w76PN37jnOfVOS3
2RBkwaUoz1LoLxJYn0OFYGp+akL3ITJSwvP3lOEvQFNAAaOuyuzAQt1+bjZbj8qAgMYAGRdS0NeQ
prx3jAH9oo4H6CN3HFm/ubHbwq3rLAOqXTsaBx8R2gOKzBOBdXBvYniQ5Fun9hP4Le8RdTQuOUJL
c/kJhwU8w0LZLR1tLp2feVP74I24G3tbnLNjUeB7knqdcyQT4xi2AUvvYifAVyjXtPfy1FlWlo/m
p3F8OO/YxDhupyve6V2sjy+STn4/wWrJ0UlLznxPhUzxM0B0553GcGPZVvminOZIEPE8Er2snJfq
ZjWkjVR3qKqfUcaV+rLc7pJivLzZ5zgLdCR62P4ke3f94wcVmCgkBK3EX/O15I1mcggrtd5uT+cQ
5SOTrKHR7UVrwgexSrJqRDSIWwkbHHgDN+ToHjCyleep5R9ZqMFoHVML+qDLM7mcyUznPUbS0nx4
hDElfuZ7+MYtstU1RrCROYJjgC9B5zMrZ6EbYTMe4/Pwi8//ypuj8DlUcpDw7uWh/uoIrtq9PhhL
q4MArJ9vMvWwXQmS6m5627X0HIfCx4ErjyXceCJUtAjcFnnoLJ49oaiUXjr+Mpb8bLCEM8RfdU+1
DA37iQ9tor5XW3nMkd24Pf3lUQlsBe0/QYJcSovVPlfNj5iKGRod+XgsFaCgqMURNAjSajPzVnPU
YsHh6QzFFHapwu2v4r/uAa7ozUbWokkFySV//LNzz3N1G/Aiys51IfiEPl2nuqh5NVP0Y1A0pI2n
d4buAfmXilasRBa6b7h3unmrOFZ4zkYbjEGPWNGp799PJBRB7ulm0fHu9kCafs2Tk4B0idshXlEX
4KKOyVTRKsxKUs4voTpW/dlglpWGsv4IHhUlxje6LlwNSVAvrkiGFW+o38ILrLqxGGrw4vo+bv5n
CjLOjdMKWB8Q02PZZSpOM6EE8K94k1RBys7kVOoaUckSjldomwpfFGmSlvozE2zN5I2e1hwm7vsk
CEZGVCFc1yiRHmwMoqBExBif9w3Z/g/Uw23QjrbUiKd0Hbt47ML8PdLCe6mnO1hmUxXWDSfLe45Z
0DhIR4B5thlTRVCXC7pTXq8PTyXZVkj4lZFbMtnA7H4XLWCH5Q9MbH3tHQZb7469j2cHlZDgcu9/
6XOdYUMVxqrTzrol/MCcFG78Udv2Cc/D4plt9rZptkwOIH7VNEwsJWwkKbfSMCXdoo5DrrH3C7ZZ
pliK/cLPzGj8odeu2T/jQme85WeIUHOvop6iamZJ8hBxoqBFj3RgMI9lZ6rpWFu+aY9VGm/zIBTZ
r50WSz9bEa7rqbb6vCERXSPxPuxS6wPfkKWkF8IqAwqOuQX5CtYSG5gmH/RNsa7JqdwjArNUB4z0
GRNW4xPRylSL5WxPxHkStSrCoROJqSNJkgPu1O1FyLU72jhXxzwfF2qq+4VDEFgHE0P/grhg7meK
pWFor4QoKSQ4V47GlT+1r1jz397MIDaXsmFvNJE2iDckPrfFN7enkayW7c1t/mGV11bJxt5efkVY
gTzTF5lrXztG3gQBYC72vExDXTY8d2nsUKJYQBFUD8H0khdJAt+GPyu16ppjkhuRmQYw1I9s+3do
TsHSZAjlm4X4NII9vCQEMGRkSbVnQR0jBexyV8ds5fibfd1WssUBdNeNSIkidTjFN93VQYDxlR0r
CeU/vfckf9sVgIM0bcHTYlM0WeyB1fL2wlr5tvRI7FnqnDRISiydT04I5ZnK5c9g84zJtF+QHIB/
B55Ei0AJ6H3fSowuwv8V7UyyqvvNCJceQY5Vpfjv1rr7cDFDy4b+DWPChImr+faxZOG1/dN6OK3/
f9tTKbuQ3DTKmy7xtwhEjQbvN7b2mZP/dGNGIXKlie6LIyhsK36Z7V7z5m/oICL9d4Jw2SNVHFBP
Z5G8CKPe17WVE0xamvNFy1Cxh2QMIEaVipcEi1mP5S7/zyEC1qKiuDZ3M/yRz1eB9heW9dJ/Z1DA
RjY4TfmCvYh0hmEz7SVB4lfW6EAv5NakJg3/Nwkr6Z62SJ8tbLRtwD5iw0hmHhDd8DqOEtP4Ds22
uoNzfbdDoCBESo3N9Ft4no/LTFmrk3SD3I6nxGLJXw6vNxxspahfgJjspkN8x0a0qa/usdwZa8Dk
BnIaRnz4XfPwaQnJNrNcbs5tw5D3CNDwZs630bCGn3tVu8aRqsVWPakiGLwgqViowMNB5quSovA/
yBxKFCpYcxo9zhuesLkoanQzMxlqeXUw8UFrLQAjfSBucO4NAgTasu+AB5qykb6j6kGVEB5TGWq4
jVNA/lqb77wQJ2l/HIWT7/zNQZOE2h8K1PwmvkcjmxQJFdXHKFhNG/5/QEt7Np8mPAYpk/Y7fLN+
FeS70KUIei+k1io+COgrEKysrY00x3UNh6MpYZg/afDT2JQ+PPBmtLGblciS6bR3gObiFIeNQwdH
ih18Ea8SpdZ8rFiUg1N5Vt3T37lpSdolYCVtky/Jk2LxjqL82qm0LJTf5uCBjBeDpl7quuIHHuLt
La7Zg9TRqlUZJO5Om3Vz5Zk7y4C3IWWiOWntNgaX5T3tRWVgm+AKd8LzoWHC2G2TPnerjQMT5u+z
t3j4I1XzTuYQ3mRp1a9ohga6coIX4JBSH7gDdQy2EQCAUVuqFSbQW3kXjszyPc9Om9YAi0EtWYFD
DFECrH0jjNM4v7fhzoYsdOD/2TgV9J8rvl5Ovz23laWbo4fsZF32RUyNOgg3QWb+G7ZvDdmxWiRo
YaaVs2oC8ERmGKFEUuvuiFfG9uXtdZZ2RhvFzssumZCB9oxdz7dHrxEyAynWjbBiAJqlSbfPKLfR
6RIrDp8QWYIcZb6u04F4V5GilkU6zSmyzzMbSLzYUS7eJUxaFOxf8XVD6s2kBdN+vnFKr/N4vGOg
nNUjBGo6LCvfYn232wYeaOxQuMOovdIl4akDDjtVpkcV6jWQ6WbM4Lo1OR4lICXHPW7V8xVH2fel
qZ89ubqlbo84usr2gK0BdByfhm/Yf9o=
`pragma protect end_protected

