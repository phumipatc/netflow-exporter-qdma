// (c) Copyright 2017, 2023 Advanced Micro Devices, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of AMD and is protected under U.S. and international copyright
// and other intellectual property laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// AMD, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) AMD shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or AMD had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// AMD products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of AMD products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
////////////////////////////////////////////////////////////
//
//
//       Owner:          cmcnally         
//       Description:
//
//          Check parameters of CUE for correctness.
//
//////////////////////////////////////////////////////////////////////////////


// VCS coverage off
`ifndef SYNTHESIS
`ifndef SYNTH

   initial
   begin: CheckParams

      // Key Width
      check_key_width : assert((KEY_WIDTH >= MIN_KEY_WIDTH) && (KEY_WIDTH <= MAX_KEY_WIDTH)) else
            $fatal(1, "### ERROR: KEY_WIDTH should be between %3d and %3d - currently %3d", MIN_KEY_WIDTH, MAX_KEY_WIDTH, KEY_WIDTH); 

      // Response Width
      check_resp_width : assert((RESPONSE_WIDTH >= MIN_RESP_WIDTH) && (RESPONSE_WIDTH <= MAX_RESP_WIDTH)) else
            $fatal(1, "### ERROR: RESPONSE_WIDTH should be between %3d and %3d - currently %3d", MIN_RESP_WIDTH, MAX_RESP_WIDTH, RESPONSE_WIDTH); 


   end

`endif
`endif
// VCS coverage on

