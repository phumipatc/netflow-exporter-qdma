`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
biodOlSbU/qDqU+C9iFC7F2uC4VHNcBFR+G/Ryw5Zec2+WU3E+tg9uWASDZ3wNK8tKzxbxPkG4fE
NBrhHq3i+RZqdqpIC+4I0MuGqgVdhzJ7Uz0Vh2VonrbLU7tTclRxpzzO/4cviQov0gMDGfZWUUHN
1AZY100FsYe3DdZYuBfiNfxU6GXDTC3GAPossavQlTTK6pGUf4/h2LwnKwwwF7JiUbUCsQOhvXsn
V48GK20IyESpfbuEbeDnpis1YJVtb4uFtpUxFScZU46fNhInhlX6fwk9OWTIcqPcBD9TF8l8vDXc
N1F0BYrc1xFLDZeCuFM0o2gUtd37+cwSu9MNeg==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
t/4NH/ShxCA4XzF/rn4aeYC0b9ZKYQw5HGPj90Wt7du0VGE0qFYk52xB2YWLR36x4EuoIvna8MZj
wnj09j9S1WjPf0wAaxSqYKy52JPAsSsUr/jXSZRWVfbulHmTwCSwbpl59lRJZJLvo2cBqFiFyzOy
Fa8/408lfAsP+CygDMopJIC+KvEfdjiLi9+kF+Iy88F22bH1nlTpZyTV4dhO+QDizzh+Akax9Da+
IizJIgrmHQ6p7Yir40JSZE+HfztLHnmnB1dLsFlg9L0qJCJW/jr2Z7+h6mUvkYezhD26CP3Dq516
O57hhnPDHTcyQdrHi0MdQYlU5J6rJ/lxTeRpCgAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
fkE9hYtNQPFlSjRK1fI/tPFtYAEt4NwbRg9E5F6+zGDw5eXUl/pxv7mj+1JzEjFei/SuxVcP2mQi
SZKiJHQgpw==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
iEoPjyayAsahm8QTHFEvP47eEpM4upYnIzc4kvUcORQprAzaXb1uLZ1rznQqsbuHESOc41GQrgqb
YK1K3wueH7Ax9QI1VyMfwppqBUJt7Xx3Xtc0bAxv57FxBbLRFtK1UdcXn8ybXBR6WrD8UYCM33S3
Xt9E+puP4vDqLWEU1FN/TKJi6QjF0MtJlUsjinRZC5jH54tbX/BvNKTAA8oLUHzepQsHt3hfnG2C
vMBQ4WSogvvkGvUQ0yeTlDjeZfWXYC1hSGKTAT3mUO5ewaPC4yMV347q2L6XXgNttfk+WcCjn1zX
c3NnjDdb1JexbsnNlJUUQm3rnSmYzNMiZ7Fppg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kdqpT1YHkNyjH64UG8gSlyjjkV5VKikFcdxjVfxSCUht2KGpDOwFgqKzIFS1Mc4a5w7i9CZ7d7+n
KQEug6OJXphK/1r1oYAUYm2cDD78VgwMbVEHDEzEsYRPSanNx8fCFLiibGsqB9LGLJh1yE+6XmfZ
ehAxyd9JuMVBQZABqeO0cMrhOXnD5M903czPEqfScS2ZkAEs+PYeWYPJUTiiDNRtmaVCdGLZpU0r
G/l/yh5dt6RYFf1hSRwghZtpqe30+OVOEiTGB9/e+j6qjB9C6hN3a9Z5jOchNiTCmmy6kS1d7dfA
ViMl7t1wZk9JEImtfVs7W2p0jc4OXXcqQCywmQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ucMh33ZcEgZD0KDrmB8nsVfwlGEAkAWdT0yPotOrvW+cyZvYtMsO8AVZG0wKVDAP3Q4n7rdmmy5I
AEwMczsTEGdQRNQmggMHmF0Qqo/+1b1Fwrlez9okCQfkud+S6lYG2BC0hFFr+NzStLdOlfGpFnNj
SEr2DIkE21KNe16n23c=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
FUDim2CKVJbTVPcF5FTlAG5MCesQ9mSEzy/G6CkhUVQ4xBZD+fzapA44j1M2Nu54uZIGNUFQMZy4
Jn0+RrbI2bCpXDKIs4dd6oGZMqelWWOA29HXW6LDCItcZjb0CQqm86VyB8J1Ah0wn9q0QWXxxe4L
Sdx5ajtHdfyJfW2X838+hXxGo7TnYF4W0B/1sa61xQZzlXsDUf823p2qPW7f0fK03it/vQ6MxZiK
4rnhe74iwE2L1Vp2LKKzGJs4Dqy2bH6mR1osHgZdGa8/ZThIZXNllcqH2Gd0x0bQ7JGMSkjYNJ21
//cu2y0rxYO4fvHGOLOQ5y9JsSrX4whI4ubfow==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
DBZn4hg7W89MsKujhLUEeNJ/EED+x4SXoQrNViFMmNZB9oqNqJb02SLsYC3tEdKIM7HcrShlp6nb
5WrKrTuQSXd95mIf2TGRKv4Ivln3aZnp1/gHy3t+5Jr76uUhrQ61KIMF3XPa3OZ5Z1hh8pvI+MK+
E/ZPU7hqrYgdaLNoOVHhT6KnZkwKEtUXCtvVBhKftjotqi+SmC6XjB5o+hUnL8OpBIwnWt+hbanW
Q+nSpTl+8BeY+Fiws7d2wSH5H35igvuHUzmU9Y2nwEiR8MaSnv7ORjGJyTl/9/OallOkPjejQmP3
EEMkx2YH7mX2MWAWycw5J5KHayNQWT/ykJzjUw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
VEJO8q6vlC8p3xF3zOPsfV52GoleSnooHeYO4tZfCtXo329jqeKr2tyq5s9KGPABYIChmSdOny5D
jJbDdIw+L1Kw1uXywUV7EVPlo0izVeTXZBuc87uXlIIs/9Ql2YPiU2bomUaUup1AoiPse2mWhOWa
4AQ5rSTthGPa71I2HVw=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
DWDSttcU9cokPDkEVnrOYeQIiCsrQzPKqQxjANwaYxS1/uzMtaavLtPXclc+k+OkOR7leWdKhTGF
+ojnHAHXhWV8kteAhE7QZRX6mcWpJOdmRChhPlWuKP1mfIxAsixcAw2kMG2SqorteS2LPEslFjNA
xll+BqKsCe+V5wmBlLD3CB6bVLMkO4+QU9EJJwid8Bfgo7wHgrXm+jaZPQ+4EZlSfdfgkN81r2Wq
F5Q7wHumVMW/jtOHBcZzS7C3CJj5zXfn6kpJxM1mxLEQP36hPPlZIGpYi8oaYEAdfZqZNt82AVBq
wB0ZHAVCXCwZVRUdznIf5q4nGL1FbDvvnbPLhg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2784)
`pragma protect data_block
CCVMEyNXg3v86EztlFld9ihRqKmdJqQy3GLwgI3y85Xctxjywgf6oEILlbU3c958H0CHNn4K2iXk
cv/w0hENqW7EM2hqi1RgwT8zwmBPwiLuzBO6KMWKy2LaImwS5G4slLzJxn0t7PJblmIC3AkaqznF
9lZjLoxoY7CpTal03Ft6iWY5Y8eS3fW1IQLAqPSIfd9HD3kbWYWD6m2BQo8B1gUKDiaUNykTpdJD
JSQgU6BFRnv7qpXP5S3q4+jLzPLmqBNeLf/QTSCS8UbhYxyDO4HeGLiRYkQM5Iw9jooCYTkp70S5
dxA9mjFHI7BdW8xYhCpt+3gn9yzPD7Hr3iocsupfbirNTIcA6j5suLYWmbsuPQozEDeY9M889QGv
KPrt2JE3SObCYxsQ9qLC6EPOEDM2S87o946GTKPZ05HI/8f59GZC+V9dLzxMC6gG0L/52mDxnVZA
gMllb8HeOkp/9CsuEG5bbHTV33QHW47TNj1/NLsjgDpxt9regP9gzasbpwWfai/Rki+KDs/vTyZH
gIRmwLCsK98oyyYYsVxOlYorL8AgNeB103Xvvj1ZcZfErYcXJaK6oroJWHvQ7koaFQKUooaO8WGJ
qDc62eCbIvHS0a5S7xxqcbGh9gVyHOgg3pthKdhrOMquYvnd/EcGwiZW2Nul8uy2ejvUOyMYNuQP
tUeNVvTEAiw8F0U6otL4BWIWxYsxCbVNHv/XW2vAm0b/rpbhv4FHnuSbSgrWu08FoK89fle+Yn5F
Tx4kia2kU8E5Ok7V3jXvTinhFHS6+fZCt3zElQ/VaZgnRoMulZoAk8LZGowUFVPNH+5qW5uwDK4A
G73FqWXc2uh4c2WS9OBb1GMp47FrY4lOlpmMoWbcjf9A51InKlZ+np0yqsO5gjZRCPA839u8XEQq
oe0BGQtW7viN0E7mURhyxvuwmbOv6WKxYshFwWZ5TGAWNwb5+cykShaTUZEXrG6cILX8ozU68Duh
bWfqTvHAogOGSoDlAOSLMacY9QPWZi2H9J+tWMav5g81Qw8m7iEQxHkSknG8Ogj6C+CwBZnZKfK5
hYDbKN/cKG3yasx4+ata2pofKE2H9urxHhXM0GJHJbsXPD74v77a+J+P3G7Dgo4gv8IimC3mktzn
hlaegQBBTJS9nriWMGM+mioM+PXfZZuqRoh3YNYYT9OVwMHkqmmt7C5x/Ioip3wkGiXTPdrOJ64V
mazBwC7JoQjLHCDHcWT0KyMljslbg1GSgeMEViS9hALQTSU5sZrUZcVsJaGTcwnGMxmrnQhNMG7w
C1AvKtausBSM1sZSf/WtclX3Yo79A4uvqDKehBDwKTqhn0JyNWpimfB/JWOXVL/gF1ici+JGSXo1
urrrXvQ5VhBSBjTwte8HYWwATYcsfXC7nd9HwmwjZF9yrnRzkcfAUjW2QzX33h8nBJ/lYyJ3sJoW
4tV/bpzonV3kbA49Q8l4voi6KQEqFVtAFMghUO5652XL9b1ubtCwqm5d5gT8OR48EToqmp4XRl/8
0hMZKtgTTRCrQh+NdkINzWHRQ7hSl2R4+RAmjAQt8IfGdBwInpFx6FHiwHxC1EgM2N/dDYuvk5Mb
NXp7rR7EVrNfb74ZKz7nVVa/ft/ueQri8YQuQD6xz9xQMLZ67yNNg7/QETaCwMI0E5KS+crFipfg
mfXXJGI9PsCyYJUvwWaxKpw9Zy7kei9hwzLAdwRRgfryX3OXPFfC6vW9vs161ZpzoK9IX3ejRGax
pQz8/lrbsmS53RJfFRb6ARQRHVtnD7l+wpOrrl1h0sBqnxI6/qOEpbZCH55xAAD92gDjZm+tgmN/
T+FXR4nFG358G8a3cCmgv+j1Fd161gF2dxDwY8kXoySRq/Icj5OpsvCIpWhUR35DwihcHL8KQ88M
WbLXhhYqnSdW5VwNvn+XrU2viT7F7E4PmSeVQF8GqVv4xPQkd9LAkqXYgpsm0zCfOqjsRl1Ra7xQ
BAiBB1NQ3GULUJ9klFPA9wJXo3Se1Rvzx4NhzYAN5SHg0yeTsm+XmKsQNfn2hGUICQZLipo3s+sN
VBTJsC9aaKmpfOXpxb23H9RmEq6wGNvc9S1ec0DH442i70oQblOBTHHLb0mohAqQEonifESjH7YN
ov83M+Fs06/AjChpZnfpYzR4roW693uXkPv+9M+oeYscBPIdM5v1cFRx64Z/ZLIDC7OE/ScilsF3
O8PEFQ6/Iy2zYaKDUJjrsxGjXf4Jx3T0UOlqSnCOHNo2LQtQq85K7rTZXwG6JAHYmxZbdc2KN4hG
ZOEplHYvZxk9RzHIN6Hv2K9Galzw+cEONQblD4tkWvwCOtTVSdusd5NOIUboBq7H7yImRNSY64lo
Qq068wBy4xRwdnczvvcqxgGcAz135LrHRAw+nqWQMImSmYLfRxS19PYV80ihhI9Wg8gqJVcAnHVs
KBRP/nvEtCCKrw5bIBMHJL7C0EWAUF5KhC9Z+JSxdrI7bDGo90C3kME/BNKsu9+uBKkC6Wj3dFYu
3sZU2azpU08vtE0XAx0rmCWCDAAnZ+Jj3eyKB0IRkVV6a8Itpo9Lka7uuExBqtWThifUwjDVZwnI
92VOgD0F7U+mfcmLRauQLo/RtFbBSXDudOoPGOEDg25wOfwlnASfbueSBrRVUMJfhh1NG28rNmmW
7RjoFW2AVKbFjZCLEvtorhK8Gw8Bw+ffee6VkVH/Q6Qt/+6GRGtMG7nRiv/5HDk1K7olbG0RX7zA
wimrV3GhA3RhZnb3Zr3FONfw0DW8ewAYpDCLkV3z9/vLYGd8uIvKRmhVj5IiQgHyLIMFmJWSos2b
VLv7uOdRizG6A4Kdc1yu6WUfcce6Zcmheo2xfxHjLJuyZLkU3jl0rG71jDm6AZ+5B5RpvzIbQXQV
L7NADcbGDq92z+SdKPr3SzkOBS72TnE1iVqEb2FTUq9lYr/GdWrVWssBckRjeDp9DzM9FnlEJ+mf
IFBh3JZV5YnVJru6p21wmHghtCxYxYcVYMe9cUAm47xgOybrQNEjqMRZW4wymUuDZj9NA3yOJyi7
S3lggjsIwmuy3jCvHmXZpU+SwSfpz38R5haFkEvN+lhEHh4X06rN7f03jUPm306eScRp/b4LLd0c
SGDQar/RqrgXeair1xgCuiqYrDILJf17Ar/E7/L3sWOxnu8KOxBWDeHrvIG2dRIU9XaVwlqP31U2
Cs56YeAXcz66zP4THRSHyNa+hWhVAyWC9mo4hTx3C/sjejnPOWKmbOXQwK/OZai1OxIZW5+m3ZIa
utzv4k4K2FuIBL7We+IhIx5+2EKuRz0Op0V2OQQQyLdwl0WlzbH7HWu76w7yibcCy2WATtPLf3d1
LX3wAkAq6ETuIVE/46Is7WrBMCY1L3yj9ICnGzPKEovrhOki+Df+q/iS2MrLGQ2nHChCJEiVQNz5
Z+m/JzMIGur28wlB0sM0QwwnJTfkTK8npgte05zFL7+k1qKUr1NCbPhE415gWIVBR6iZVHF9B6s5
yfdA7xDFl9ifBjzlScIHHEzMS3MgJ8PZFFPlCZ3rUTTIEF7opnqkKxoXIHzd66SijK17SZ92XPUp
VURnKBXiEJ0UTsxHLWHbjVhU3hRCbL3PfGG6Uogr+TvTYkljurFzsBSJs+BZg65tdwku/4hadx9c
3kOWy735+8ciaiLc7BpppZ4UOU2XKZJOJo+50uBTUuj2dpkr8bDA4ubOujzB8tOe
`pragma protect end_protected

