`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gjZ0QZRrztDtxBJnXheegk50kutU2qk40U+BQ9CxBgKw3ZBfc60QbERyVeKERGIcZIXy3VCDycQY
xzhXHhAwE461BTS7aZS+dBHkWbIIXNg+Hkcy/Fpz9aGngxA+G2VxxFHAX12ZQJn/0BI9rVeSONfk
SkOI5oBbsFfnbga0cfEM6Zn2XQZAWlCD3CS4THfeXEWmLNQHO2+Fqe0tv6qf8t19/UCnUDVsZI0B
CEDRTdYjiWsYnYoX8XHEi3PaV6pbbZ7D5qUVuJaSAFnLXfQSO6oRsphvFPLydaB/8iPbRbG62NN+
+jmplbXwEw9IjOpDTjBzo/yVadH3qO0RtIHYeA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
MeaYcFkL5Q66A6Ud4sGS+LdLRu2TMA4tv7rEX+yMAQBpfkgYCFxpu7/xvf6BLyAAXO8Zcv71wstA
Sc1s7NZGjVWp/goBuxfIDEHQVfckNJzemFAYVU8P6JuviLszH/qOhUHliWVvEjYWJE0M1pHtBRwV
KRjKoxvrkAIvBcVya4RaaaCFy/gjcCdYFrt0azD5R0Zf9ztmVDqf5dxQwKczUZnub9p21dvW9//X
hgv4j41M24GpcO+sfR5sKUUUv3mIaHcavnewRz4tbmCXuuxlKoofmV4KIRHleT7zLFoRN+D7Dq9L
hldCkYlEniatEklfMX0XA7PT76Hx/wmPl1XtvgAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hzN7CSkss5sOo+1S0Xr7S2WT30OX89Q1wKx/3GLVQp2knVGd9X5RafWjhyHkc/ihs4EAOst8FJQt
pHctrgRKiw==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XvCCSOJKu4vLN7USQ3sFQh1BMSzWK28D0TSKG2Q38VqdBc5lJUoBl5KuUNa0eJjR5oWPM0zuDF2R
iCrmjV8pR1UgUkrndrsvqcEG4NBxg4JZ6pCljX+Xv9lz+pz87wug6L96S49wJ0QmCJKAqVIYMe3v
eqnwxCJCyl4PTgytXSeM8TyaJv7HDUV6F9mdPj2VS8yQeoGK7D5qTvOT+hnNw7aqDqp4S/rmSD1w
dTBaMJ37LZrZoQKLJwJPybVGxtkVhTvn7DMrYqOQqGVJG8r57aULeulnZIKROxqNzAYnM9eZvJG1
Xrmij+u0uCJmYla2bOGRsd/8835crEPHw6pRGA==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WGHswkIktju8awP4N+uFORu6on7/0X+W6kNUfkW8/KhsRGDNVw3LeDn7fMLrvbuHdrmmEh63k8UX
fLjnRK2lfVXuHETuDH6LWbP084A9/NYRZWUdk01kNv+kYoNXGWhY6ZkUoOK4sRUyFOzXn4R67K/T
tvv/BIswbwjE/8/tla49JlsFMYRa9Tv8kF11AShA7StMuIoW+vVc1nz9oab0nRox5xwUGo9kLJjv
Ddnmk14/gNHxrNHgkvwYyIXg/Je9yfbrXHNTWxvV3ARTlnD+DaQgWuZo4Q7KwhRPTgqFDPYeZaCw
iOGrGGhZ8ozaIy6jTwFLswGGSBuquvDhZlKksQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
EvVoM0fSrj8Oh+IY+kCNWhRQI8QG80nvMowXgO36e4/WLraJaSGW3EX4z0EznE2ubNOMCDyqSAcN
LrgUk87aXRO2OzzXi/RIdcMOAnYow2y0z87Jrg2HT3Aw8FENi1+Vf7rO3NIO5Rb3GHG64NaDOhjr
Hx+B7LYojN2dNB1QZfM=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qyNHAnbIeSSojh3YWD6BjQHaVpgQMkC427s4Ax05QNxtHF51Dpc+iXyMdakXQes/oCHnYT6zbCJb
KccNmYBw8SJMd9AOmTIn8DHyZqY99/ES5ftywBKcBLG8vUk72CG5Vtgw21exAVZYAwoQesAv0Z15
xJC7MhcqCdlOokp49kxpGlzwlXxEeftW/SyJZ7C6rqzza3qnnTps+b5R7brgMBKRen23lelbtagp
pkpYpKFCJIYRPlXODCLGYVM7Kd4dauNxim9CmEggOEucSU4nNvcjmQKrdIELChq47EC9kVI6ySBQ
JloA89XYsSmMsJwg319Ql8WwWfxShxcpFOQ6hA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
pfGQWmz6h0y3xg2CbdiKCdkajwSmBZ5ZxHNGA6aM9d+0qEHZ/ffYKgQXisHgUTz5emrDK4laMiVU
4CgAd5HRd7dw+89VvF3U5kISlT28fkOQ03u2csajAD8On578qReJlhCtEGezr1Ds3ZsvmhFor+DH
9SODsS2P27nOVwChQAaC9N3XWFKzKe1/dUb0krA1dL8GrHru0C9exA6dK75HbIpIc2Ov6w8oKc0Y
ZmwguVsioQ1RHucvLwoRu5kkia6bD1AdipmeYaFuP2mDp/oJFr8GunFaoF7kmcn3B42r6ENJXulS
H1Vuqa4uy3ArZ0JVmT2G/OPMHy7E+Bx1oavQdQ==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PUvt5iwAgtP3KP6aFiMNz6lY7ABXR07SAqWj3OBYdmcAFOfk+xys4rTaOJaBGhxuR4iJZdNofh+m
JZtc2psmjcriwlPepPmg9IlCV1nlziDRJeDdZp4hCGlhXVGutDOx/cKBQ8NMZAF5Yef206mXxkED
wYyMkWDspxjdOYK51vU=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OXITrs9Al1GDDI6/9dkbPpR4hmoS5p+lFHELQTSlbuTfwc5oPrUDIoaQhAeEdelbAIn0PwY2os1+
x9rKQuOK7wcyT0ShaEsTgc11bziVRzXJY5baKTPLh47k5PDivv2Lm+iLPTkqCE0kcZjoi0YmYT03
KcgUqA+2Pa10f0UpuqVzugJWqvLQ0jmm3UhUaJdhnJR9yvJ/b3L6hX2agXntkWGnt7xrnbxoMvB2
KEhZ7/HSLCgVpu23rq/k/jGuzN/RcMb1ih2JOhR3kJiKF30kSaYZtX4bqUWSr4ybeaz2aOYOAMfV
jHcDnz+9G1E1UVvi+cuyrRETGstNjLdNOmztzg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25856)
`pragma protect data_block
KQDWCGf9uIJOwgAoAXp2wKWyxeflhWGGdHOk4DbHxQHlipZ4LHA3RYvbagBep0KAFRBJpQiUusNN
mobHCIRQndA24FXtWdgWY+5E/2cJmo6ARPmR75xkZ4kL5ElyIIO+yi1MuD0ADeMyi3WMABUZiDNx
gx/WlV0E3aaE3s6Tszl4cXIOenw4z5zRhPhzOZZXqJH9Dna2W6670lomVD/fenVrTJUjOrKdxmUh
LeKaJUNt3L61VIDT562tQz0zo++kQNfc6YJ504O8BuSOq7tcnzXqaAbiGB/hbuQGzystkiZt4g41
BbGxuD2yo6GH63Z0bQh5CwpMCS1RgP0V2EC65qrLuoiNhRUSKDBITpH/L4xLecj7hrWp0JnrEBUz
YwWkWdO4vXyYCtw+ArGJY/pn+d+f1y8+K8+Vu25T/976wiPQhZyerk+Rknh3NehkaOZAOELsiYHb
ItR/47/O6hOULOzQLXgp1mlWszA8rmh4CrjxwTsuosl2JK6eevaMppFmRFoxKuyfvDFtoTPtXadT
zDfMIXvRQVx2IDRA+z7VuofDb6r1j2bQaHoIPWn5vyPVfuOUkgOM1bim3pN1VZImB+GNNF+3VeXY
tlPQ7SliJbRuiuqPvC9jlOPKsWNFfqBvqWw9Ay4M5ycY/qX3PgKQyGH/d5UN25fqfxJZ8uf3Ewxz
eHiepQAarmZk8b0udqNp08fDgX7BV8FBjK8shc1MUZwI3LJtzwqmjhJijrV0G8jDBHj31fnFPxcH
4kYceQMyRik8Kp/VlTu6SXx8GEvmwjuHqlZ8E9KGD2MqDKaNC4OR2WP4mXd6i0suJ1jQN3jjoj/r
7VOcWdsDz2sOUeovKlLTmZO3QF0f+KDfCvrVm1Uk8BwtNGpEDc/rMzE3qYbCDr1lJ4EfWtuUvbsh
nbQcxApEyiyMQiLxXTWSqZTmAdF8NpxTrDqbFjxfuih3hFF6vJkDF6oQ1M8Aib1GscD8p9BMcBHv
RZbbUEtw+o2Fg/3192o0A4K8VhWHSyGoYpe2SinkJGAvu2vz0R0O01gKgRIjvxV8tnSpuuJB3HvC
2mwVUQtGbYfYcED8IZq20KVbOa7E7YqycyWyksKAr6r4rVJFeovZoBNfOp697CniI3T9i5sm8Md7
bQAI244XyyCsBCj0NIIrWhDYsnCBkeCj4lRfZBvUQHXstEs9BrdXqAAcWTMZfaiKi6BDrzXTh9Ok
PgPt29dXLd7KMXSn+CLFUllPnJNTw7QRPJdFoyVPMsk3bzXlzB7QUFpdF30lZoUiKCxo/IuJ14aP
byVUMOe8XwlVVP/+nDLeuzpwuiODFlW7tjhVyVjizWtQfDWTrJhDvyT1s5oJQCKgVaco4B8VT1j+
F/ay7cTc/9rtgkAO+DpEr6FW46oy+Puwn/4Clhwg8SGklB2ToYAJOKRrWLr9t8RyQon4HqBk6eKk
+KplDci9QNmQkZWyELj27W/5pjIub2hlmBrd/GkIcTdO7zTqJ6iZT8AC7LHIaZo1936IKdn4Jnd4
ihlYTniCaKyaDjEicL5mUo4rz2a1c+rcBDK/T/ckqq04yEMJNXSadln72T+Fwb2f/TPUiFijWFXM
qBdJ+OAUUOc0Jt4j+nE1l11wpUG+EDNkk1o7jWwS8QDx8VMbO1uNiZvgPwOzkstxFjGnHZ8c+CeZ
VbrBdzV1Rdx9pZW2Rt29QcoGZSWU53AHZ0K8zogTDiirEv/a5gYoFqpjPDAVFb0cEnaKVnUnnHY3
w2FTvX7NXAys2vmw95mJBgUE4A2yF7MTl37Nj4cxB7mHvVLf0yFIG8C8YaxlUSg5KY3yDupBE5WW
xg4uP/4D7gRnhHi0EHnSgty0mOsAAeaF8dgiMhM+YGC9Aw2hxd1RYJX/HYLheDJ57sZP56RtjjAK
yOMZfNaO9qJQLJGZD94bxwrj5QEqFET5jcK9pC4zL2KFP44RRcugYDIz2y6Ha4qSTgQJEEH6kd7M
rdWFR2jTxYsOs+Cnlq22x2rxEZHP8wXWCk+GeKoh6oV/ZAqlbhdp+dwivpkMpLSEsoEu0Yk3Z6oM
Uin3VoLQuraBIvSgxdatCBnNRs+neIUyNHFGKdUmecnMu3Hs4SBATq54sAnw78zA/OVVuMyprLal
ehaKbccSDJcQYp1eyfztaeaxucAD6LMuBZa0XBzPR6gXHcHTUWRlXfdSuSckWC+ChURcBhlr7DDq
m85Z6lChpcE1qFQ0dJHq2rMlZbfsQPS7F4G2ojQBuQ/twD+nmQtIOMec9I6m71NlxUUxsYzx3MJp
c+64wPAeBB8720yRI7SettvNsOWATFvpqTp6j/SG/C11E/7lCXyFN74GmfUcNlKenEh0DrMVPaLm
PCp0lLA02kv7HakZHLs6fyxbmMzF8xgg4lRTGebgmCYui0MPc0Ie/+PyiZ7wVcztxCb2IYjTctvA
uF541pHs7HEAwIjkd+golRwMcFMrOiZNHvCzSIKkN7X7df53wcRbPX8N6zgIrf2uTbQ5T+KsC/Mr
qpG0NgG/OS7jefV1FHo6yLY3elFjwzxwEQF+aSWFORt8K/0Ny4nL76J692LBaJUtoy27UcexFh2G
KzIUrbNAMEKN1XW4bo5j/kNNZuViEAzTWF9sbRtQjVmA6j32Znc5SGGepbErW2GqQgQ+l8f5Ltmb
kkpItO2Q/wfyBL7Cqlmfv/w4vhwV/jWCPfmXoDDukbIoLKOJKDIRMqPUVjYoecUfJIn0LaSUs/Ll
rwpesfIupgGwNQkTBRYaLOtX7UeRYBU/y99Sd0uteR+7MZ6t7jXNuZKKH35e9emovqSUvTyeNZyt
M1/QSX36EmVf839E1CAS9dtEeAYWBXbD36rJoxe7zJqmYpONUmLwqEPAzueg2ZSVfxreZagKCcxr
nk3EOZXmYmzs51QVeuRLq1IkjUO8DIBDRymg7GPy+6XWLeJw4JG0yDp0TmACmka0M6Por/BYOfF0
YNZZQ38gU5bxzOpzknmUrr9r6XCkrucFwBp294ttEsnUuGitQOXFdzRc7efJ19SJehr+IYwGFq9H
Np/Th4jpbR7UScIgBdw/h6dDReLdC8ANHSrF9YzUCj9lo7uB/w6LO3lBNZVsb6Ry1AHtttVceBah
lYFh+p4VDD9PpaPjB7kAwosWyA/iKyLgFhZVqBUFjKOCN9+02MbCsTZwRrDJIEvS+XNodiJwpfJS
b72+gPJp91FT7nse7WBAEeWuChhLxXumhYwkqHS+oOYu9qpDeVxV5fmZKkRC9Z0ebR0l36lcna21
+VeJQSo/kD9+BMRDcPCCDWgSRTgMelqPwtSAX7OzTuSegR5badAhAt3TCrhTNZez0ljGzajtA6HQ
KI+v5W8kT1baUJDahwGW9QiiMLbYg4+cl+ujGQPBKX/PXqmC5dMGC1T7fYJvsF2uij9SbJ+RgTY/
Y2k8fYHoKkdXNPz9fVPzQTdp1QWLMUQWzL6a9beYyCeZQ98rslNNdxcklVLw3I8Hc4IgGudn7E97
jLovH8NA2CSBz/9BayVcSGincKef7h/iPVWpgm4eR/Uhw2cU6T42GIn9RuTPq8SV+O58LOQ5JdyG
LQJDNWUHpD0OnY4zzyXQX5B0YrRQBlNTDC4a8e3bYthNZgNd6rYj0xVk+chu4emhCOgCuKk6ilqT
5E5zgf/HReqpCFsG1gCGrLqayGoyNFeybTSJOmyWkVFHD1dtoS4p2VIPJJzy1LOnJ9Ahgl9MiONK
YhKffoXw3HxU3ss1KEKKi0a9eol1C4Udw8a/VvQTcXEfL3fFedQbCwrYO3xmpffFjbCSsrjzjJip
XnJFr/nXk/DJfEzSAwgZD4avIiAalF13Gut1w3dNPioqhR6+GwqHA4QQY6bDZuPj+LIim7TnM85B
ZFIKPHGmMuG/Ii8Y+ZEOlEsrgU5bmZvUmunt1mqAmSz+wcuyacFxqL+E6JlHHmlcUtLu/Q3d+HHv
yTdZoyzI+rw2QS6btgKIy7QUti+7iHtqePRrXeV08EyCBEoTGabt6H4Prfd9eO3Ja6ytcSe0YX0Z
KeYNl8CY2kfi+zqNBQ3wWhV4ONxOSVPime+exI+QHpgSi+h29O4rocA+PEwMN/eFzChvhgLh5u1e
66e9sNKNYTYf33OEoxjEA1jXQRBSIQqyi7bPHymI4wbmsp7KDUiaZ4UfVEx3qh9UvEvm6BEPk+eW
DPtPIJqZc5qU8WSczdqGrEAPu8MzRiAueKSV2/7xGZFOpvDxw11iP7QsXk3gvNyCbUYXgsBDMF/G
dY/NpoEghByiOpPP9ONdMjcupfnfWhP4OtvryK4zt5gbYllY0xa6Q0LH51zde3a4UTtFSwzgNOr2
zrM/kOtlM9qgRkBbh8u1wd5oVV2ODxt0MfNErHLu3Cla4k8JwqqGYMJAgPkcezhYER9Yj+59ME0I
8lDRCTE76P+rkDqj0bL2iRvv3bFYRtJHfjtLwgxb3WapjDLv9x16pOqR5Sx1xer2dO4jdXKQfLt/
LFDUcNr9LLjXB9FqFz95AeI4avhR1+VpOKvFIO6wzvcG5u8zD/Fq1942p0/ciVd5A/eQJw7+2WWL
P0/2xkRCeifFzqHPIMJtmsjn1O1wkEP3oP0m7eYkaHJSkGS1QGF0hbUiytFJAmt0aTG1gWhRdOy+
wsKmnjADXbybNztgx4Ad4jMn89HK1b6CQ1gf1RwGEJhRNot6riC3MK++q84CNG7T22ECtNmSS7VJ
fhf6fmdHNei1dDG6mPB0JEZ0kHt56dji2roLFQ07aF1GuVi3/xAqCxq3Ik+gWrcixzAGlXYKaXdt
d19HOfZbubILGQxnWGfN0r4C7E0R0xYQDgro0V0331GVV9/ERugo+XP/Iiu4KJCrF2UmlNMIGu6g
FLDyy78H3F8UKkGo15xP0mdzULt7W71DfDXJLTKGOdwOv+EdL5EeyvaJ08vNlio3chQOTbCyk0yO
abzKbCNdYfNbqDTGiE6Fi/fhZ1VH1ddzS3Jw/LNugTN5nYOnBF3Q5w5RKok6bnbV1tCsF4AfaLln
UjujHbBmmnTCGxl5U6kO7PZMwEkhjBB9th8LzrPTKxtmelkRB50d+hQxPY/+gS7YTgCP5POuI+T4
8Df3K20YEYsYoGmoYUKq65oa300FuqxyjMynxo7+9ywHRqKrp6v2y191z5MEP2XOoDvALEppeD6k
MamtnWazJ1xyv0mFiKCW3IfnjjNvwRE5+0RvNCGSLHp9HyCFH2o5UIj5AIL+WoILUPTVykN+OBfb
RzFgkc2S52FlOwzAOAanbJz2c8ASbPhrXuwusWE82pbpDyWzppobCw/S32yySKRFHfCIZo/Fj+MF
2VcVZFWApT+IfKCmPjUR+GDluMVoXF8uQkSL1l9rZVY+nv1dv7ExjHDSzsglZaGangokVXccMp+j
K/bzBR6xZWhy3lF/3pyekEmGNEcFtbxHYvGX+shVHrozVJjBFAwRkPGcTB25k63KSQmirrsFLg8o
vBnd8SMZCQm5iET3RruO/xDlAvWp0FFskDosWCMmos743ENnrHyGs+uXhVvxwRoPDjIqm6DnxyAU
Gc1k3rre+GZQm7SLeCTh6e7e3b5XyKtXPGB6BE0f9nu761ph6tLA4h5JyA2ckqE+NFzNfBUvQDqi
TqQKZwzyUslKpbOY6FC6vO9ggcbuOyaZ88SjVVaU1c7nmaxf2CpoTmDi2vEmiKBaBS5W0c/3ctG6
ak38llF41rKKWVeaQNcDMDHi+Zfzv/5Vr20TNZfz7nnHn7pqSDya/FmJQgSzn+W0+yxPkf9O33FP
Xwqr3cVZWK66x44LV6l65oTmrzbjPB8J4PWRv7N1ZripDII9t09Z/F3G3+/+MmIIX6Wa098jDVk7
55UzWkAGX9iangsK4kXUU+ouCXgmhxA6XqoJoLvzIfNU+DrUun89mSM3oluc2tBVekZosaujABL6
NauB3XcAgZWrgHhhO2v/Nnko3RfyB5H0Es2H6RSTXNk/EVydnhVpxoEy5St1t1wlXq5eCQMeRAQd
QetSuejtTE4tBdJ4dVAMALZQGJID5kNOtFzsSMFD21nzyvuW6Qds5njxzj3ddAi6yu+gG84wLaK8
uUpkf2Ys9+RlwWqaBEio5XSRSXU68QAXaNC8pcFxF2z/ddUIrFq/pzLcPZcQIFjiwKDC3zwtJewv
A5Ze7bMZzsNC40hqRLSy5jFQCeLFmssKbkQlI1rF8ADBfOhnJ30a8WdvTlCmVtLls1bdL+CPiLCg
wVAEwjzYcHLuJPBQlRRFTSuABO0Ua0SePio/OpWwleZGh2hxHc6/zp0gj+clVS/r0eZqNkdVABlX
C7yHlOS62TNZ0921XoIgJbXPg2oZVMscrOGAkd3TiWNOKgrHqjtiXFtWq1qu9h590Pn8Its34HWh
frufAekjNVoiAzNqq3sWcK6lp8yCZNr8/IaMif/qC6zLAjzLu8PT3hYG1XkgvuRK5nuo7pCyXZQR
OwchSF/8vzfPURkKIoKYtKckXTEkbT1OLbp86ygNbNdpjmj4+nf1yNRi5nRcb//e2vupGZ2ECM6J
eEiFmxKiQBg1GX1x6jjNStS/TfzstRP/WF8nG582fDl8ewaMmxeHYjDzAqbEd19undIXWMhJANNu
KvKoCaD4AXLyNQ84o+Q9UH4R3hvz6oSNUb0aYC/IXaDl7UL8gosVME881tSLhYCN+mQ+B+x08c2W
MJ6KVCR+CcyIHDtP5QYy2tKzffz6F/Wv2WpEG7dSh48bZWwBinb3qxmw38dMsjY3YHNE0ixe5t4a
D06caUh05oyQviAH001XU09614/qu+rr5GoOiiDSQ5xOkt09Lplv1F24oP48MZpr50WM78Phh4gr
JN6brGUOAljm3YA+ys/+unJWfJHiGCtcXgy90ZGbheObHAAOEVcuxQyqz+8LFlciSsu12eqzuEIl
ONELdbCwfQQ4TymUnBO/90zXoqdWyxHPLg+q7zRiJRmuTkG/giiBl/p0sHZL6vN6VYK8gcAt/gpC
u7nQO1KxsA9OBaCNfuXObATs58iDzGDCsI1dOVGPgNXUjQ0lmSjah5k061BWwxxZ3DFUvmb09GvE
54Z0V/fvN7FWeVLYf3YHO9p6p/uzAa3jSyzdzYZyAUn3GLD5RpirsdiMFTMvECZj2zT+rHJns9nJ
NUZrqheBu8gDdybiVFhvAHL9DnZW2A2x0oKbUrlCidef1SQbsAv+QTEa1DR/EMYFy0xLM0LbXBP9
1S9I87MJnC+eT0I8mSH7ITNlLX/PAFUqDQ+s2r+q1l4AiSrDIn1aRMo3UPK9N81U06t8n7zlvDM5
rme2u6JrGusLWw1Rnf/9os18kJSq6fCLFBIFTQtyR9jycuY6IjNMbH3t4USfWRMR0Y7/vLyKbEPB
fmDoyX8lyjfLCn9TQ/oooptbmtGUwNssWL8RY4iN5rbCZiRytFkXEXgyFNWS+6KmCuHIddMzSyBk
XQCSg2JS7JWI5TJzbR2HqGXTFado/dqw5YaBAU6p9gVvdmCuVSIEWdsYXlBdfPZFxEscEdgOzD9E
cYHs+Q+aw/jGi/Xg+02RDUsPmy7wavvRy7Rb43CenjLaF9XhN7U3lpaRtvVHOuGzibmWt/whN0go
ngfMYAF09cdEq8cMzSHFl7G8j5t9hO1YYFuLdyiRoIFeZISa2qEUQVxG5U19EDSPtveACmUQJvMf
RU39wfRWRrpGRBDDiH46PCcxoip4pLKQ666X8ivuFhYYN0lAZHN2dBISklJPMHc2I3c9x5fa8fze
CYQj6FcrRold6vJN36U8+p3Ip0lcNP7vrkG3CZzE9EPjs/e0/+VeCkAQFpF+J1yi4FaF+GWRZXkC
0sA9/DLtH91Xz20ql6iiNn5cqF8iyNMArgz1LdFUGm1AJAjS5SNGISQVXlT9Jvd6iOyz7t9uIAFe
fdOYhI6IRLjUHYtp8ZbZUQE2NSMPh/YsSJCCB9Wu7Neh9yA5RCHoOCkJorRogjuqRce31Godh6BU
ocnN12tIY/DW3PUYn7Gpl3hPededqlpXrPHi76Hl+wv8KxmZB9+qdHyK2erGFsC9oUvyZ4YJKrQJ
kUIzhIkOQ7zbBNK4skIs1kfLwYfRtwWPoltchcyGfJ4nYSJPzEU7+kihH7MWzw1ftCh1rg0w54ch
0LzeDh6xX8TormGv/ODNbvqvSr3B+plJRn4itXW0jE2zQstFxfF46kpH1x+H97PXK8trCye/aaLE
qV2h/RII0XbWcJfsfcfzHYGkKquyg3xjbOMblpQRZJCYCxc6SuJRe3ucqNoXrqdUKAg0i9dF6CoE
LZE+9tswNdsPJZFdTmMm7JKUf4uj5TmLOkntE8ltD6KvNbPVVCEyxhmc2CZ8GfRF9L+3cNTBvStE
kxHupe0QS9tKpYn8+BnSaSDHEfLizaBNxV9SCOmWzp7VHzYCts+d3aOJNHWqyd6EIPEA9ToYeR7I
DTfbWIyeg8HbAQX3X7FKTQPea7zi1A0zLQ4xzC2F6Km3/W+f1mKn5aW4l014n6zvJKDud/cx+kOE
UEQyUoOv8OlLtgpayADm6w6TtN/oj/vn5mZ/GacgaBd8geG4I78BeDzPisDM2V75UEMlVT5dBOEn
RqWhjNwSwKPwc71W674ZXUy0bQKrjM7qbbjIGPNA1ykuv9usJR3oYi5JI7JaW8HSIqyy1SOCz6bE
tvWYP8SQ8h0D2Sne0THMMe6QZ6TKAa70t0Qlvp5JM6m4CZd4RA3llmaXqAfqGtDM9aAUZv9b9we9
KZcsBpBPJfmRGdy6zvg0AgesSagdvyh3K/sbwrDafUbKnOv9qkwhQD8xWsyN268XL3lVaBLG6IKt
AtNXpe1nDz1eVakpzC9MtksGzdACi/3Iy6UxFUjtL01HR/lcp6fHwpdFEhzh6TKrloWT61bYMYtR
Q7VHH6eSaXOrWjgGcY2DaK1+4eMMnV0fZ1EfMYqWgFsg+e4qYs/ogM5d5GgvqPpEBHmwD/jgT/1u
PsrCQ2yPv9hlMTmRjrZgv3/vC6ZJVBoMtzSdd6tHaYrWyGDbw+vG3JZzgQfi52iP5CuhzyimQUtL
MzTAMYSJGDRkm4OwoiAfTwZXm38qdKqHz+fTv8mToLhmqprZI8MvTqsRKFBtdW5Aae85RTtBI12x
Ix3Dm1yHNVz0ap+awKED6RpJGMBNk1qShHK1GoiLalDU3U7pBQ+dyYJ/03gh2auZ89ovZeNstqx3
0kyoaH6swCcIojdbYG2jOXC/2rov1uekn7cDf5fcX5A1EmKwn9ujUvi9BDgaB31YQbdC1vA2rfJV
RskTjD6RBG8CwvqJBAbVUTTM5u4vyC/RaGWzMUuFsENWrr625VfxHWOvuNX2AUJh/xH66RQoTdRN
GRY+q+Mxts80UOnmcCQUEiZVShvUKgjLAKxdd0hCQdyHg8XAUMnoHkHlnVPwFh37CH/8k+QzBU1y
Cz9reeAdMObNhi1YODlF+1PaBd6svnN/g0IpBSoRoWK2qbtWILirxg5wEKfNQIe4rv+zGXBx/VnE
0qQe82WBX+2mXzWTK+wsFfAqnDNYhtkXfsJRVAwNBUUN2kQW4b9WcsHGRDliRKKWBQlEueTQFfMq
MbN0I4rgXIFkue8Hm4WKTZ4lZmseIuiHQMC5Bk3et1c2Qw1tWtXcpvCQDOcT/UGd+B+xgjszETG8
oLxwZ0ByL1UoSWebXVDt0k409jUnpNuFSjehBD3bNO8e8T05nIe1ceHP72nxmQpnxS0PSsBrL8vf
96NPbyy1mZqEwX/l1ZLjPL+pPvV/1J3e1C+S837imnI5WFY4VZUQVPCGgnGkS5qdAJjnApKcSfai
4qykidhEAf1HG46mTGLoru09X2sSx2ABaOm8gyl12iOF58HhwR9e8/Wgrw7F8SqZkScSgR+AvB+1
PzTrkVw5gYw4cndf3/25lDrbCDqG31Q98WXhnMxf3fnfBbbfGdXdH08A3j30YqruAzcYGpA2KcNP
PjSY/GqBAB+Ldbm8pofHCtvw2lFp7sDVxLDaPUeAh6kKrRARi60sO+4ktkKwnCagGzGLUCargWAe
jQHpkm1W0FWqNf0sfwWuDdPBd9eryAeLiHtuIe0C6JsjF0pn2Aq/ZtHPy/QWOiS0e/DIPZRx4lJq
CtwSdo6xioEvK4njxF4SHqebqm8bvyyeLdw7wud6nWvkQWRcqwH88isoJphZsbnAR628iJOHQHcK
MYpA0rK/NpWsxQBgQviaRiuxufDberaROw1O6B9LyZcUSpSD3lIX/Sghkmaw19uBh00BE7pFDJqz
jkzV5V4fxi8r2AlbVGP3wPk2KLfiIvmw7oC9nLhx6MJ2Rq+3wkmh2cpyu6mk2O2SNQ4c3e3ezwR5
5ahcmJJ+FQ+EfdezEbSEduVz5KbvxwiTjuvjJCiLTgx4N5nyNLtLHa+XwqcuFhZ5rgYTi1+zY2tH
DhG35fT/8N22Ix9o8H3TVPySqUBCN1vumSbhO3q8jo3Eo87FH/JU+VedfMrR+VFXDKVizBniWhbI
lKPjRNKbUqzin7d/B/1ubgbhuL7xhS5gPK3Yy0ZPG4OF6OsOeBG3MDIAeKyxYVGlxyVi52c1HzYN
BrKj/bpO0KeH1WoZJcswXKIKBB8NH9oaxKW+8i7R/euC8Ijb/GBIKzrm5IzfIrfn11TqlkozE8sA
g+1tsXcNfUwUvEt0cNjavctEsWZQ4zIEIfW8s0qeLRFD2/QBCyCbT9jMFX13ca0Ku4wyNJt0EsqJ
egCAruXDQCv/4NVATz6Y0GVNTpNmSj2t+9im+q0UIP8kW2oHjglVbEXdpXg57GJsro6ZE7J4h1kx
wwO/q1I63fmhEM4tNmeYOToalfeAhtlEeu7lhawa5uXQPfiWoRJ3yuXBG3hFMEIIxDbAxjwdIz0q
c9hmpoIbVcR08oujVGVS/s8tsTxCyBeLa720peEo80xy4mtFwBovUClIed0C9OlQrv5I1htE/jzF
WFym+xBgeA5Hs+KQ102UriFhy3zGzzQetZgqeO2ptetOAHiTP1Pd3WA6RdNfOMd2hTSsWrmrE1SU
/PIvr711xx/vUHucJXSdiihDZ+gPVmzocfnp7wJjxn1O0m/rCOti9FEeyV2gtZVodROa7SyVOasx
me8X1ssKFcQBdIXTIzFp+UyYn3AtRcm07+LOzZv4NCfTsaYXpiFndMh13miXkyQ555PPOrAzGEgo
oNFsnb9OopqeC822MfQbPBbsuxRmA0ivqw712xXB4BFLOdDb7sVGYlDgnyt6MCI6vpChEg3LgzMR
K+NnWOW9RCxw7ZcNnG8NRaE3E9664NXVCIXAmDks1OhttBk52z7cL4NtiGgKiqNhz6pvkrcFSrL6
ldYzJ6b4HtJ/dxXic500z+PxOcyVeQpPGPYVOtuRaqexpno2wJXnD86CArny9nbOwUALmLNEUCwa
6whYGxOVrRKAJLgWFxN3bvnj/P3noNmEvUH7RCdHj6t6zUUnT4d+87+4VQXIg9gSs58jef4VDwJE
FkQom49curkp8bCs20A1+U3M7NOUHmSPAZJfSwFxVkg6Dgzoe8OFkcKFuuFrIkjfm0SJtpgb+vvN
3vuixPqQyXVq1glQpnqqgSBX9oLeLiRr2JrA0O7VcTxdDvJMuEoygBGZNkxGK1GNbv4E1utI5xcG
yA/Xci7YiXceZPh1JN8LRxYW6M5cxMKEHf6K3JuEfm3VMfNOwamNwW7kVg/Ex8+o9LCF/VUIMKLk
OmU7TdUaODOIvE5TvIc21dzGfug9vAQvzjsNQI2T3iGkzU+fsP3ZYu7K71tYn1iDCMqxyuVgYsuS
zUeCvw/F5KcPf3yJY1erlMuf2TcOQdsTNH+5KvrCkNUOWFzZUR7l8RgOj/c/UPCJ3+jenqg0IJG5
s18jQEGKIJB0mRdnhGeBWXNrbajtbhqdZSgE/vEFIra/t8D2v3G94TOOg+cLZRyc9yu+CWrFHTU1
LQ1fRluMss6AquYeoX1QjBEJb5m42kAQ3fTbif6JMX9D8yYcwb8bFgIn+D/brGAgErVgyW6dPXbd
1/MfNu65e1h+1gvS8ZVIUOZZEVaD0dCnEmS/PxJf0W+EAObWCCNnQpYHx3zQhDE+uPFXaOZDFLgJ
j03TmusEC+qW/lOU93+IFLO8+Wt3nwREBsjMbKSkx4KNuz3dhWyhsAjq99EnGv2OiB0AKB1a2oIn
2lzCKqYjVpv3srAqGA29G1Imf0r7jMm5V3V80LtDl2b1Tum2xYlDxvshI88Eqd2rKg1Rsao4HN3d
If2VWY4uwVx4WgTDjmo9F4byU6/gxGKDlTmvME/pk4IPMCwxE/grftaJNiTB2IT8QKbc9HF1Sel4
YwjZ2JPeAGWuM1OYDFeIWXpWHZ5GlkNsXoAUGeUPhMyZX4iRwJ78hkqSBVa4tcYK8D/ufd0y9smP
GE6V1g/ZfhK0umzcQjsOYPAqT6m6K7Jav5RJVDdWSsxzh7Dz8emW5LpEvJFUhuqhbAgYwEbgxDFr
rA4/5lot27Wf/fgmnTB1zuMa4DTiXHoyXSYEcFHzQSB/iHTHODxJKAv0Ixi+HIOUzRpnle/MaxvA
i6+3+lR6w/M4pq+siPZlvEmp6sJlWrp5lesW5Tmp5xYADXIulYVZ2y9d2rKptwJMFVgEEm/8ZQPZ
OLUGCunZRuy5frPUPCl1/UtXOA5RhwYwrbGEHKMi+9ghyQmThWm1AG7UEjLlk8BvTrTT7FF6dWXS
L+WofOsxJoX7Q40IRHwMh2ICrK7H3A4TKlLOqPHeGovQJ5zX6zcvwijiGcqM3AJdYYsu2TvTnX1U
YurXReTWyNULxZayhWm9q7TCBmAotHH3H9JCWgMHyerhfu30QkOUJJn7ShEQkaW7IXuEwuStB2Ta
ZaM4yGZmLRMHTInzo4j4CvBRQrBQH/OdXDrNpk7/yH0ey1NeXeWKwktIHPLev2Ddi61Xtkk5xDUu
DloODaxALA34UqQB+eOw/rGgt2xKdnJeJiQcYlmkEfFf6EDO7l873oNOtIw0jFf09cfcgN0ZAKHc
avGax3tF/zYLOwE3aPgJoh1aaCBVvD8iKNZ6znxcsu4JneDyHNnbpONVW6YLsle27NR/8DyQh+zb
4Jc4vUJU6gsDCwBXHTYWa7IxHnAGUBj7T+ZzWRJOb75nxfWgrh2UXGgMK+BmdfRq758HPatkZ9wZ
VLvDOZW6muJAGatPAohhnPc9BVcxu6dlkZFJTLDJrSJmeECQdbXOEakanL3bNVwRwhU7U8LdgTyV
Tr4rO3GTUqLcwD4mSiUXCHpHQjjnWv4sQscnU/KkTRKTrI0u7WMpm6wu+K7QGHom3uAJMltw5k9O
RSb05P2VEV1n9sXKKwD1Rl/E3UkcKO/OyEJxPdMh3G2Ss0HecqBsSL4yTOu98EBhSWMzMOCG6Ibs
ohYeAdx4A+/GPxzkES7RRkW8AJy1koKO1pIoq/aU6OBwQVP8qXdh0pQkAZDqJg+lhOqqv4VQ3yuy
jkXPpJMrWLymv46DHI5oZmeU7l9BWIgruyvzbuPGgnYVWZpvrY6pSwxwrSICdSaX/K4R/1s/TTM3
0nQw/xG/zwQw0TmuV0FrethiosxQDBkT0tn2031lAlw4LegDjPXtGnKXbBjpOm5loq2b5d94wks5
NbccWCM+4lVGucNOoIkc7jzY9QECwnBJcqOkc6LBOjIh3eJE27KA32Mc3fO7j7aZYTQgOMvcfRpz
8B++TeEsZ/V1NC6jQ7Efkd/mNNFqnbSRhEPIn9bLX9gtUcmEtkGqY9LGXWy9kokyYO6eCMcDMY5H
5VXvcOcpCysXEgdu84tDrrpiHWkxtrGaf9k/CpyzPFHyVCWNcYqERf/5uYORkTQaXuBZ7XplVwqe
dAGedvqjRAMb6i4tXFgJ/rI+Uq/TA0DA+i5FXq2Tn1cGBIoR6ILFYZeA82vUacS5PMrqFNRnFNvu
eylQXOO2tbJYQcdlAtv8URhLP4Dx0d2b9uN1uMRTJidcpda2CkAgSddT5jEvOOvxzh52HwT6Z+G+
EM8aTOxXtQHAovfxp4DFhkQaV0XgrxuGzj6h7ibQ/0V6788OpsLdvislOF+6eA1i7XtFqnBFuc8S
BXPGcREaKbphTCSufgI8pVSWfFgU1nCyWR6Tg5UGWbKvA9Zv+tn92YKDelCuorDNQBYvoYWzIZmL
iAB+yJk7McaVUSWI2DRh0Vz2AGcMeY/0VTF2ioao6J0lLePYNrQJlpW5FM7qmM9FA2Sjgngq0JAd
m3Sc0Sob6avnH8zbJelaLED4fO26cmTGXXNlxlhPK6fslx9ys7UWmW+vGnVwnet33VMJCXr5mHP4
lisxTL920BVyjDK3iUV8WaFQXsquZI/M4sdRhGda9oC2+LCIoSZKicYtIshSCdhVuJTGnGG7iHj9
XCrQl62Y24Kmjm23KyQLJ0KYvmAoSATnQW99ySLknGEXps/Kv9O06UCoAGCaYTo/8MGZiLpap5yT
9EyLzJPbAUwKR/QK4ya3DOs+m4xqaKjqKRahY1Q/OwJlbSLbVEzysMOYBH7hX5QgDI/QyH3Nrf2Q
JX3GldRF6pfN2dEwyyE0RaUT+7m9ZbI+/H5bbdqO5zK0ofjoGc7etu6MvG0pSEglzo/m/iT1QE4x
PSmxrusfvNaZ6heD3wooY8rhDhQgDxvASlW5DiKGkQDWuY3Jdf35Yq3o8YcQBDUSsxXUILiA/CCr
4KhOdPEpgIibaNq9yobtOW2w5fjill6l97G+H6BWcOWvfgKXhNehGkjRlfOTUXnMrz+S0s6xBIJB
a39wOpDo3DfVTmGaPRf8moXl5N8LWB9FjoGrtehyD3Lls3E8QHiSDaRs2rvqakjUrAuw7K3e/ckP
ReJGHJO4Yd0yBkN0+Mj7/rAxc+SL5LNHgR56ffjzmGpALgduIUMiIOWH+9w0wdo554jHaGX7vPnn
F2eXgrM+rLsuhiy/OFQB/u/LFLy3utq2puYtWrJSfGLK202B1O8slaU5aAKG9VH+TH9dbHr9XWob
YzOM0cAcbLW+cSjeGdEqjyRulsvce5Dq3XoljfmvyEsP52EIq1DHAC2Sph1FSLHSrhfv02wQFG5k
AqjUceSWTQYPu4zXyasBp9JEtir21XPnecwjnPbOq935IUJmOdeupn1tft/LTQgh6BwWJwBGUkth
pWffp278z74Mm0WXGl9FCiLzOCPntOBPhdXtlh6bF5P0tWRg/R0+eJ9nrrRSR6y/iAv1G7ovNs0G
34qH3zrG2YlK35TgYPMaj1XOJNKxg3c4F8t0Z7jV7klOqoY2ZhWUYdPz8QYAfk6lhXIG8B3TH0g1
GlWI/BVWMOS5rgEkcNo9TL/WjjPs5SBbv1dJuTtypV147A0/nrWvwfScZ04VEO2gnNxKmBWt9Kt7
GBY1V6H7mReMlZ2dgwlGYAHcq9WBHi1u21Udr/fmevZa4g9jB0ZdCL7YAOLDcszyBc510LkjejEK
PqdMmMLtoACd6ze/wtiSwvl7esUTOVYtrUMpBGFpxe6UPpgLVlRwqtbPnRgPcfLNRUymgHZ2C1kM
jh0q3cRNONUryCLZgis5XAzIgWvP7/n4f/fSy682EX3k4v5+bLxwAYflpRDQeRNIBjG5F5vDisd1
46NXuNFJJkk/V2ZPrGd2nceXZmmWiLxCM+lmKuUiz0d9ImAAg/3oAbPsZqnGNbsNA7tPdzpS8Hec
D2jHGoUgodCjPF47DkUfQY/kHxDXH4sXv6VkgDPkGjepZ/Dyjpk6UDotzvLaVAXLsjmBhMxYNza2
eaZ1bigpO6yux8dV87d6YfoSJPZaZRos9JBF45SdiV+qKwusPthU5gc3ioM2zF8ljguIW2PVU+Ow
SMlC6tBC4qtSic/1omiGLWbXo6QgKX14BbKMNGO5x8UT+H/EGEtopF+2iQgczxYNFPix/8Bnc/YW
2JpxtuTjiK8bqgviynezOUBkM+myJzLD+yRUkgt4qqYNuDGBbB77A218K+p+tpuO8At1Zgj8xrGe
3hdOp5urJUScZxhwoVBSE7bEflmkjvIYMqEZ51qS0zxNwKNDNl3yhluizipHsrmvoXeZQfGJdwZB
NSFFIoRzVm+DZ9ujtQYTZCDLbTcL6Ditx94LjJgRUhvlJGf3zKf6zuGb5uUhy9SfmA0j8uWZcghz
0NfA6QaJAM2mDOMfpZmSH2k8jMnjxHfVy8p2UQTrJetrp9UC3lCCIFrwBCWEHdOQWe2OYqvbczxL
2/683pLKoDXoWrD/qwd2jr4lfRbOlc3UqQ39RvuWQt+FyWjSWKkGryk3KBoYiNUbat2keghYc6V2
tEUSbMS7v1Xu5oin6jFvbsfko24y3ajZclbqUUPO3YtVNBH+lnVeBxEP21Ww5gVoiueWJVMfW4kt
0597sq/k+7kcP3s5l43x4rg+jzGHEyiRYnUaGmVtN32mLqLWSgi6TuB850XmBDVLpaV0qJmHg7Bd
OIN52j4po6yTCfIqxB8F5t+8IVjCygnkuJ9MZoa1CpvP41TTybOqIzurRFilUyXJxs5Au6pJTadO
IE+Uv5vsffFUgJJX5KIwOTXsfXgOMuh0HdZ7FgB8VLBP8TP/+XgWf9fwoBArxw6OR2gFop9nWUWb
QFPPLIc/wDfOllR9AZNrc/CQYj1tKLiSbWQdarJkxkm/BBr6yeNJWP2EqrHWxdYyHsyBhhuxSyQ7
uPt+9klFT7f5kNBPRIty/K4g3+d0hf9T1Sicxf+MloZkzlB9U/nABLuKqvCZJ4Cl+rpes5ZOiViA
8aeBtdQbXqiDZi/CNXVzUPEY7vZMA5MIdw6Pl4cIjRs6gEjwITSUZB5qaikukBP+1cHXuT1CLYr5
xFFvZzPf93jb89HBB6UWop49dAu/iCAfX95a4YWDLTWWsdlEw92PR5OprUonNBxK5z7j5rYaA+Pl
TKeDmst6doyzLzrBxJRRu3ywgz212wHYAZvJ4cEWO89pZY89BtmRx8D++8rXmhtggPsDswpeJPp6
/ii52KtSZc9j8LLtwW/4iJYwcxHhJLxCdCL+mzrzI54cgZdK3jEkNEa6M7pppyHBhmq40XkUQxO7
NU10p04WYJcbSJP4N3MSBM+jxZjBj4Tc7CymrdyNx1nOYfuujisGAoTCbdNuuCJvbc9qUcq2Hqk4
vLd5uOcbck7LNNmxqxrzGRe0olK6kqVocJl8hLb0VlDiedWWej0lM75GivqNfQEHEkwrB45dMA9z
KzX0jyV+iJpGIi8ipzZTflptQ+aTyFb4K9soBSbiqiYnqieEQtWV+7xUCANBut7RVM9d0kzrQHuE
+vKi9BGFfAsXW66nEwxe720CDCpIKNX/VPz91cdGnZcuOLuUzMEgXH2mqRkdbz52vGO9JBhYkAtt
266ezTYMzdTK7hwc69W5y2ViXbCMYRW316T4vD0RyX8/XbnFnL46TyHSSoit1usz3Ps3rKGqT8/W
aPK304eW3DZzW8nOtP6sHqiUWS7Eckd+Wpr4F6ARHW2jwdkosVkak4RzakyIRaOgHQFoVqQCozB/
4U8ty5/XIjA5ngoK1PuAegI3Fa9yfRVk9IZ4yMJXmW0tJ+negrC77OrYzcmOSvns07v2W+74X4JG
yV0otpFkC76f+WwpAMRR5nqqJQOH3iHY9QgzakRi5t6QkowKGQd7XjZoS0Rt/jyIukOzOlNXFOLq
KM7+RT7VMudEixgGjxTC5GCrz/Sg7gbCL3lj57SkrAGe5H90yZiFyd0K6UQADQQZ9qnyGUVAISxh
zBN7OaQNK8QivRaNtE+3JkT479RCVy+hjpiSxPFZqAH7xYQIKU5cB6V1nZY/JgJP4l8L7KRLZnW8
TPwGJe+JVbEgXKoC0w9a9R/Q63KrJ/Rn5e2ZzIvyZg9TCFfY9G21fcq0Y5GLugto/zyBFCxl48Dx
Ps6OQSU3fS5u+hzSEnBwvbd9gSIqRavTpTEg3+tRMS0ItW2DeiaVZmLofVBC7siLY2Iuk8ZAUPoe
G9F0nLvsZtXYr1w+gdQ2sBxabuFc33TC4SYWf+bfx0tHhb79c4TiL1LqZ6I6UO+HfgXCWyZNolml
3D4bcr/vt1cyO3PQ9PGe5bYDFH11TwIcLAONLRumr8pqLC+9Ogzwf5cUHvMDr1MifrX1EeDx4Dv0
Zjbm/H9CbeRZR1BY21WWHGHulLws5Ot4CFasMSf6uXprp6OvdVWDKfC8/BQDVzAePKXrNi5qAF6V
3SpprFd6zm951F/Ayi6VgcXag8v+a0zrOo0K4dusvOr24GVizRKlkk6nzB8lvPIL4dH3CwwjfIqO
/20qOoUVKloXOwziT8yQVw4XrowFjY+n5F/vLzEOeOMHE81Q6KslUu5cMSPVRb4pevwh+TyWUSxG
ApmMGlXtaNdVtekAJmrgZnMedE+e4aUbVpnepCdAbi2rbYQ8G5+5E7pKqRy5XtnpcLNqotQVeWrz
XZr6lRNwQOllrP8TB58r1XQPfVrnbcmi5/zGxS/HO+/WTT9hDmyF9+fKspB3Eja1FH6Co8UK0MPS
dTdYupXh26fjcOVN8WBepT2OD37mAOATGnk7YdD9ai55XIaPOmYjXWv/+t1mqrwjWqZu5pbbz9UP
LLyY8j6xVgJVZwjsjqggurVwxx9gCju/T4P5uJHkbp/6grxMSMKIwuZfEB2fUFWReMlkpb41wkls
PH073Y+/RJbw7dug+/h6UBxVteoAjTyXBp1+ci5F9uclzsmVRjgB/noMB/kbznbAM6jrLfA3KfOj
x5SNEeJ/aODx/YAcQ1whGtrzA29AlxwpCSIaFxWTHpIk8Sjf8mty25EDoss+qnHdBmmbb8t6pHkv
xlbNwQI00jjiQG8qG83+V0XKnzfrD+ZorM5EbjNO3jNZLehJpsVGXQw9KmMxRreZCtkmF50Sr3px
P3rXXGv6bTLvuAS7tOxA4FMIQEDe2OezrmpsL3mAYVsEK0rB0rW3q1VQpPq6YOaZbdsaKWSTF5j+
IYVlM095iDHZQPTX+FWcmTaPaDY1kq+10/eOXHUhdIuPhggrtMFavnYIDv2mjrGbxSiAzy86th9x
UGu79A4YSUcSp8HgFYqKoMfGe16PlGE2LsHElVEXJXWfu86g1xzAoGwoGRVi5eZrBMP62r62xptQ
AXbNwiNIUFi7DDDIA6y2z1FbdFKBuCHjulLBumfAa/UlNsbmS/cjD0VVLMjnl7aoLRkM1QOKojYF
npx+HYIfIS4MF1CQi47PpBzoGebeBiMTDIIGIUl2Zq4pzE7a+Q9lABtpzW3oMShqpg0aVg14AWLO
WGsccS2gf/bvPxUYJ2xTaxWXxFnZupt9Xm46zfkJim7uPcr2+4RL7oqlhwBBTOHDUb3KtnPKzqRB
2An1Ldtjz9KCIrpAeqzWk1tguSj+vs/zPyWkXKhrn+rN3idxYhpfi1Dld2uxOIXApsspafHMQj0P
0pQdMM47Yoal6MEMkZa1VhDo/CT1IETSWzozk2lx7BHqaqtQGy0qtwmgSSde1nzACkPBhejEUDH6
pzcVFoQWtSMT8o0u86jPxvpNv07APCYXuyJ6DPvc75oyw1ekLfLu1RAvafVe/snUzVEJIsOlzyIk
ZSDFuO6Qa4FUTi6VjDwTuNxKKG7Hx7h9Y16LtVyXnW0s9UVzTQCCqest2LWMxuPVy8C4EEvjnEAn
0qTpgkfsWNKuoZ2iW8SOh/Lp/U6OGnzZCr6nFqx3BB5NbZ1W7gZ5dE7R5SXtt0wTUuWyFbEH0lqS
UHIRRqFYgDPKwXTfDiBzVtIihJ13faabzSDFA48+1E5LM7uTMGypPd1NXL7vcgdkRgrRRVEzYIre
10vGAtk92EN0ar2z1tI89+hD/33dEeQ+I+LA2MOsR6UVGxU/G8Sjwfb3ezPoFwJUAMHbg23dam3Q
aPtkYOv8VTEvLyUW6QPjwzhAu4nELnkPPfHudqlqiT/SNxNGJOHrbqqrdZLJ2esNXGMt2/oN1vkc
Wj6dTcb5VfY8rMFFDOSlS/GoQ/8xGU7zQLW4wXdnBtMnrO+P7egVWkNHnDNBITvZhJATxzdFMFrL
kfq4EwgaezoOdrnbYnP6ZDJekwqI8GJAp1OpHjsNzHPIw0C4H7PPeK3/jLlzVCF9Kw2alkSbllrd
eTfpITGlAABSIWm4dVRfnicZYP8jSIviTtqKCONoNl2O3xwNabB+QEkBNf+05s0CFk0S+BLcQcpJ
cI/kaB5nZ42hMqSij5UDROx5JAbVZIFtpsfum4NgFkn4vpAmDjXQI68ewpZEId/9iuuQTElDMEbn
KmLo1RNyXxiqfxLnMxyzKAVOfhEBpckJmckq/RwTfJiR/C744wfkPvZsXAFVcD6FuWg3wQZDgozd
cjBJ8eHflr72cpHJ5C1+1fOedtLinzH7CnmrfXIKWui/MyrJZFdcuCQ2qpk2DYPswIecPhxvugZq
bTWSbibPV0/5YN4cwp3yrtu1E/f3z9q/PBdKbT+qVAbTFKRLmUGFbVvZ7HeC3qpXjRoD3hTPrvHH
h/73EG3RB/ek1tgmfFRYws+UEkSdVpDATVwm4h6Lxg3NVMRDz3PvNFMSDGAuwlz8gXIoZszPZAYA
2nlMjYd6zVGqjrD6pwHGARYCaXPasd5J8T9/cCrDnvRs836scocFcmVlO5GCxJ4ZOWSHVB9pThxp
a3pEe2GRvrzL3PZPfn0X8UBbtS9ETXYRAnsGxpOxjVJ5zSgMv2HfsedM1zUMhumzOMAOolXOK4hi
YkGojVoWUH86X1P4eUqS9YW3vSst7RYw6Y/Oj53slsXjVkz1ST5JuGbJiHF+0lG6nFyLKU55Xn7F
oxmmwSYJwXEgWl8lVNlHKYm6dEcGaRXjRPY5H3KLmKQ++5exAen4EU3NYqdrDSmv4xjrg7LEs24n
wrzQDoUnACaIrQKHMk8xopAZBaq0byVSAnBx6UZB0Fvd4/515gdug2Tfkq5axLJuStLcyeWNyAu/
yZn/jj0cPhi5lLIp8CVg4j4EEjEBqPYpggq+3T8v19Rswl73tlYAB+HNFZcLRuBddLc09ceypJ3V
goig9fOZqhcf5w+QHbpFW/2vX3Pmgtd0C/zBa7HT5GXQcbni+8NMA54mHkO/r0SeV1xw5RxJnbhF
tOY3L7OOwq7MU0hBqgGSgNDl2tF2vK2NQgom8IQCZXmJ0RyhfNoH8PWFoYBS1jEGhPyMBFnXMu2G
bvNoPoHuWoLaCMdZ5x+WfRPLHAjYjUo11FBkP+pCAGOiuDHMvT2VLggOqtiX4TbsTNcxRAbBhHTN
4nc+1nyC36DXfB5ONUBvwyx0YnbaY9lcOuhzwgsvbx/I7Lrw+CAdX7k57smdD+QRt6oQcY4gw2Iw
ii+11AMbzsZqYY7wiETTsr2SQ52LxfR+l+vns03WlAz13dEUPZbda0r9TxH4XPBoV0JVNulA4kjM
Z2+Z87j6Nj20dKbBHvwf46ykh521/wqSQQaiHnDcJk6okhiWgzK0Fp9rlW2GWYgXAjVxb6xqJT3w
0fTEbIUHLFLMTCow0dg0Inf6GL+mnKsvIa1lbuVo130IOu3ObJ7Ls6+7quVutxB2JxRcn/mek030
U75LP0aaQw0dh3toiArZ8pNV0M39/IU1bXBCwRSuP5YN3qUPonRbaywUpplPfTMML6PfzFdguCYq
gfCB6si9A9AZPWPW6z/uc1vWNP2fwW7rgWiYLDIQAjYuaSgAQP+TDnlpn0NGcSnbSMGojZi2wZ+8
RtpezPwwAVWI0tgEdFq7DmIn0zzy0h2ryXprBW9zQKFscEQRj0iZG85emndYTmEaJpEp1ggNbMZe
Gbycv0AXPAVNJOxO/xXVCtFzE/iOqSa+2M68PrBMv7sB2+EShzR9l8vKlSs0m+R2Fb6U5d6uirP1
aJAxSgy72zJMHHLjzJoGVDEMv7PemOZ0VBxAhyjARoteTf6ondR1c5TBazBkcSTVShSyiV+oqIvi
Dev+3Rt6XTZaDreISipO2F1d+Q08DBxpw39baQO4vx/Zw8tSNS4pUZzVzmwGVNZSFWgBia4LCZ+Y
jGpYOBULs2dQZ6TdBUHlEz32XC/1P7WIlTXiDXJv0Sn2U5aGto3VyJRO1fxyJHMfu3xIAjBvrqGw
PzeypZG01/T20VBWeA0ZiI7JeRpTdTc62sHB6IrrzI7JsUSfwmwqNHSpFxvWAem6xBufb0BeAvsi
5ELQrZFeo1CJGjifntLrVdWMCoPyq1tLCMAlIaqPVP1JHbz+t5eqpwaUO0lpVv6Y6LtVCnPqBipM
JDZm4gQz5ExX9xbkI3h4nhCxXuucRmY9pbmGVGDayTgXAvNAyY1enUkFDOqk6erK6bJ/YZLYLJKB
Ci5pdec1Gw0H909Wi+Btdh7V7l3dyWKMVkqNjXPJpFg9M+kmtimmQYGvXUTW/EBsiQkgRIxNv3Ij
nPLWH2KrH5qrImidFyUTad8QcO8TeT0oEfyjGXE+HV7vsOdDSacZx8iX2Z7N5Ux+AUdFCL6HE6ue
+FMLH73pt7kjX8yvPSTiGNT/MuxGu0OZ6HLBDnY9+4cyGo7weMq/u7t9YZifmRbAY1RbRcNpyMJx
f4YvudNjpHYi7O58Yso8Yzspvmk5o6jghnvAbLEcn0lyHG8cKxFiMSbMNrOGBB45LE/qFskyl8/9
TMtjy3hOmNNxcw2P2WmkGsmDMi7BOcT1c2d9Z5qZhOcyV8ZKS8jjnF38R37TRXjwEOaBQtzdeh3r
m/zVTP0xgrjRpDFPuK0JH89yOfAojl+x5VYN9pKwmQTNfzPhs4voJC0ou3XgsYWF2kfK+QLr1UML
fl018SNkwKa2pMBhMblWoM+kbdmzZUGEQjR8XiDCE2gMBlmu0vYmNBmGUJJGkmrv10if7zRwT3Q9
l7DON9EZ7KoQHAsxTtpy5gMygrOY1QMtbeNaMpl/2TwTcIl45L7kVt/NAGYABWc6GwW9rdxLJt4l
DWL9enz2XqZyW+/uCPmC6mOn7Ka2PXK1c4wqDaE6vQmNYUUj2dSVLFd2lOtlLkZetwIxJayT9yRO
KXyc/I4v/2h26jeKQ9PMcBP8mKTqX6QKgd8PWYaYeIb2esC9ChXy5zOYJxQWeVPACB8/JRZ5BrL5
Ns1ng5mS+07XS9Jc3eobFqyCNsNwdYR5gHZxvbxal/838W1f4g7T52v5Ec/T44vK6AcZMKhS4aYX
H4lwvx1GZ9HC/s8gs7Im0bQHZMNW6kEl6onA6euv6f5vCvdj64T6oIhepXAp/oBQj6jqaonFOKjC
Nac8k2FQRaK+B37qLrYJDrRhTbX8i+CtDX31lMbOFKf8PMqZu9Obw6XV4lzJvx0reQ1JOV19/cvA
Cn56bEFmz0GLh4t6bRJk32GIa/lZ5rKS1xqHPVrfrLI67h5eFLBLq+IXNWF4lG2a2CqKzJ9ny92Y
ZPA8V8s8jtPv+HpTu4r+vsU2BxJkERbpyPKMfuT7GYx33B+n7HjSQx/DUaaZax5TVYVA6dugKPak
Zny9naClkajKje869Iv/dqxfXtYGydl8VyYLxx0RSxf1T6GFPT+jmyJ8bgYDgjCqEeBSpaayggVL
9hNRqwHpuL+p5Itx5Ss/lCcxJum93g/Lg6kQV5Ul0jzB7Ht1rpYWtOU23Q9mDOhe8YkAcUP8pHi4
iNczrh9Lb57IscplYxSK0kU0MfWkzyDmL/H01os3EIdChNigwVBffp20JKxqHR6ey+u+DuewkIuL
knZKZ3HI9isdfgPIEGrh8luQOEUqm1DJah60At1ch1I1ut1SIWCkw2C4KKlxwRhjTokTv70JCQ4O
aHsDwbd0fYoaiZkH2xKJ/O8180DIUkKkNfwJebPqm0fbbJZP6WM7S17Edl0S2yNlMaHKVVusBarZ
R4umOGEJngYygBxYL05dc1cAkz0U+5o2kJSmDPgTOd2uS3TCjJ2a6gY9CknyXO76mOAuDe//ZWdS
Z5KGdv/KAeTKM7zUn3taO6105o2ACzAyRWcwM3wgnK0C4kjg4Qf8svNtnOKIzoJGNdsFBi5MHf2H
DEScujRf10nP/eCa7ONZ9jpPRcJjPVYiVZyJE600i7Cg36C0kLjNxWGVrhzPS4a1/n2NZ5MNysiO
GEPvpcw5/WCqCkU6aZRoHR6LkAFtyvlrF6ygflb971th0aXsZdArb/nP94wGqphO0fSXvkyv6n8W
lmhAD+X10J2KEHINxG/VpmCwiWA7XqzOpHUIlF7YXhws9yIdXVdkL5aKLTjTI1vRbY9a2Hbc13hd
k1HjUuNqmwWnzBvWJU3ohzQ35E2MQea3BwLp9pQXkkiMcvXd2vlifhfa957oBTsC84E1viw58MRT
mvcin4JCVQlEWM4QMysw6PDZBzH8fj0aRQvfg1UlqjJVS6Vhg9Y78aF1fvzPDJzOc8mHc4dXgW5v
GyvBVqv/gF5Y4rWCPguHD9xNSG2wALaAsNDKvu2zambD3yf4pDifATDhuxC966XHFbVgirkUxDSv
kXUBh+oWErgYmjtb1FxBrJwgzvDRKDA+5d7NmAhajDtZJJ4w9GSr+kf4mPQmuLUerAZEvtUu1NI3
uhNk3cUEKgShXCQsjOvkdvA7x8vU+4Hg5GPydk3pSHZtetJnU8TcM5SeR/D7fJEpXpXyaWmCe8XQ
856A2xX7kyI+nDOCOELb3g27aRtswMzkeyc4rIcV4zSuuiq/Q4n/uHQBxD+cyXK5MSOq6q7XnWP0
p9O8iYK37ASoSAtapCcYClDLTZqx97nsBGe/oCZFhsEYlUgG5z+HpEuRIqi7zGNBaQukA5hvGmC1
4X/dVYHZDxM2OtwSWa4bR4CfanLKujl5k0ln8OTQJy/gTDB5UOeapg16+i00Qts9MavXIHMEGBAG
T+m7L8eJCVlfU5pZVPPypzPAv5Vp671hnUoXUBB9K/PZn2tqhXgPJhd0iPYT+OXeI9vcPyuvIMEL
P8gTHmgl+pIfusf0EgAXKl8hqeKILEwsCE3ydtmkd3QZjUvGCYEdJNcX86pe6Ar6svZdnKUt7NOE
t6kfL7jHi6XQAeG5QhefmuNIPqV09YgBqBUS9GMiLIskXrQhstQ7UlxCthMHih3EtDdtnTHv3mID
UBLb9j3wbjnueS6sjK5PlZa79FbZIH0jdyk1dEIvrYapzzfbarnz0uz0u/SHDDjVdhZ5mpDy3j89
60Q+8a+i9nrq2FqhQM6mH+Ezd2WBIKjzzFvxiQd7VLFI6g5NxItQRxi+OICCVq3MWb+gakO4Xrg6
sMarggJ9G914wZdOvuMysicBeBFpTXL9K/tmQqZbU1UjL3NKFazEk10s5TvfnE6MHnk+ko+7qREM
C/55Lb2f8XWN4fXfRwqZs+A9BnA8P7OE3wQrMK6JitK95Uq7sT+/cbSkp3xL+hOwwXkd3CHFfyOH
ulMPZxtgSrl1CsPcHSED9VJROlahF83JALk5HGDIdr7ysTqPP9oYQL0Q7td9n2auGd9ykbZQuhSy
cQFrJT6KUsrP6e0wrWzQp6zyuWLbFaCkIrxLAQTEfnfbmn03yJMKRKclTGAgMmYvvI8zf5vF/vjR
U9vQHC5KrCm6aIr/zVni73+TEZmZjfAdVSRTYG5Ijson0Vie2ZgROXuHA/QaWtOyhIyfFw42ToiZ
ns2vDpka8kTu4HWZZiqCpN31+0vfWTel+2D8oWmEZD0OXgwT6EH30XbzgcDzBgmFS/dPY6OzaWGX
nsFbZFKvIipH67i17E5reDxOuTw1T7kPkgw4M5tA+PCDUIoVTUKkjzAfTOluoWEIRJ+YsZCykA2v
zICy4TEspCCrkHjNOrHLs88y4/d82Q9lAsSJlTDRNubU62Az0ivEywpbSyFHCl01mzBQEyaO5ts+
C6r+YoEmiX2OSThp7tYQNtWVmqLqzwrb3hUKE5kzaOKmGVBj+nJuhtwebK0o4+I+qA36CXW63GIz
DeQfjb3nNj+PRYUerNNqsVtzBTdUf00bcMIWueSWA2bBVgJdkrPigSrkur0dYY+GEbLRofk4ekki
CcoUGBSkHBExPLwrECaQ9qAHvDj2XbwDQQq4xnhWeGUaGanm9DqFbaxIf0ATtNKkxJNWAcwqa4GR
Ob6QfqxDyWqDSEEkRjazLzXkw/+AUurJgaslJKxqtYkvfS5mHp2MLDWDhSTKw1rEuGzc9tAc/i/S
rPmoOS6rRFWUVrO4xsXpSZM/pmfnH0P1iHO3wuoHZFGou7eawZViY6gRVU/JukLWR5SWs5TYZRx6
HbilXRYKWz+7Y3lHEqKFOMO1pqBau6rJZ7y8Hp0+LljldLHIJ7XEAlx2ki4Z2q7BKeFZ/lg9NcF5
OXpx2HU5O5x8/FdbbYWW3VGNJFAgBx/Te6wE1ixxvPm6APPJiPQ5n0OiNKuGElun29KE/WZMoHI+
3CO4dpqyXXisnh/cnLKIJjTXEEusppaTpIN1oKyfxl4Kc/fkvCHk0xWHYe4Tv2MY28bOE4C8kLzq
0bsbvY4pCEnbK2JAxRiyV8TafB2x/n5Is40hrr3RtAXKx6WWl21/ePKpmaglICWvPWShwMAptIjI
H+8zwMvTskxQdJqvnHTV1fIsGglJCjpigDU9jaqRPUtOuSNLBTzKkUPeblXxoXGNopiyUnVCAxID
OvnzWJrYSNSIFJbgcrY57OKniii8F7q79X86v9UQX93uyWF8UezsLeJh+AtNH8zPZla4H61Ztdf8
ozWzyTuyIT1jSEFCNqJ865MILo1jbU5DVtts47nCbTKQKTaFHOyPPXuUbgyHVPiD0dPYmFkxL5jv
uhHZf3jR4LLZmkOS2V/1nb80RilbcmV6L2BtJPQyMrOMc90PAVQx5ssno0qMJ5t+BsVWfOcO7Vlb
3XgYxnvd+EpJBFNFaXDHdLnhUn7JOeA0Dx+tvmAHa6aOARKc1YzvrXw1ALjAu+U96JsWd5oiXjDW
AkCLic4o3P1zXXGpqk1Rn7UiHl1GXRELQdP6b5QU/yN+BIXGzMSvPn54qkC0h+NICFtmNWcdTeQa
L1eo5pCf1t7+IhFehYmdh1FoOzX0RGGw7Tbv4N7QJHmmKzgUcA2YVVN3QUR+qv7Gr6NL60tPZK5y
FYqpZti+IJ3QITpLn+qtlCG4HQ7sp/11sDUiApHuM4jyM7O8yrvX54xuW7SEnFcih3A09IWTnCng
7gmQgRXIltrYdIXMbCKLVZFzpyPjfhT0KGOM3FC9nfh0DKfuX5BkzD+2ZdwD/4/QD4+4Ldb2dTjR
+eiXP6IZBfdZrcUvECJV4Djtl8IVD5izs3ydUfS2GV06ukOdaHYt1TNQGvF6nuHKOuayipp/p4+1
UxWI6XNRFj+dC6ZFtYOXgINC9aysTJWo9svDqD27fF7/P8nCaZo9prbMqmO26fNzZdtHXuUZpyLw
pNEDYXC4+BDg4wyH/RFBJsWeqIvCAGjXA2XHrzM4aEDelCNLh7/RGcS3cs5V92gKSg2qiuKFBa1L
9Z+VX58hZ/0Qhzq7qFETooPzRK0mzyz8jq5XsFiu+XHi/l5btpjel4pmAYwUmR3MsyMwUU6J7PCK
8JpEPAAkMn6ZMj+rAfP21HMB05myvbLkcvKR8qJe/9Jc0TUciP53dmcdWseiU6dW8URKMudZRQoi
K0EvyO9AhnuD1k6S8w8Ufifnvqq/+XjiTqS+gXGvpZC4sYBNrTzWngKCl64s25iSL6+YEsQUC+xo
dil+UJ6bIRLESk5bsyRN5owctUm3pvBxrRCfA7ZLHXAzTWj64ehMZSrddwv8NFNWalk/YizGn/7h
S6iRuTEZ9LEYWk9RQMR+U2wtf7inbNqMqNI8V/vzeQsQas+kPPv4NmVQdZd8YP5yGpw2cFdr9kp3
w9FI6gnxuTfHKdE5RmemxQJSQvDA+muDRlrrLo/1uDAe6uD7A3QFuEGIV6do3Ol4TwkFgeph2VCk
t8G4bmBvb9EUUTOqkj2K5zTHZ92JInUVWGmLe9KJ3BYc+K3sk+vN+E+g/QgHLFz6zD6P4xdDsLrW
KfRH01K9ynSx/DitlYr5FCq/8unOl6Xxx6FXKziPwtJCkaztAwBvco+sLpswvZ0lZ5iBuisO76cR
29eiJ3mfO8D71Z0pPLeZXSrGwgZSY2uj3c2y3oTpcdh891/WplWR+W5QoUoonmr05bkKqBuRJqHL
duk7tou99wnIedDcM6FE4sQtxG9ad4qMqncaWi4xj9hGFtZf9nQdKPJevsnfLqQcdiRTCvRXS8uI
kvlI9lfbT0S2a0qfAZlINiDFPfkS+aj0N7x8XqXiJm4BW0vOm4JBGgG+46JN8EO29p+IY+psUWK0
IdwnmuEESu4NA48K5o9rJVX1D8vedEYJlFhzU4/WJdycXw36L0G1qxPg915JECaodNMoEh8X25MO
qe5WTFzILB91dcLIh5I0pR4uBGbkzNx8zneTYubPd58afYF80T4HNzahULohF7iNAPfxudRNEJv6
asxBhh0+3riF47QfT4YUC18/gi8H0ZM3BCfUBzEFIyTlUgU63wx8EherKPTdE8MFMJ4G96l0VWUk
wGMIBib7fHFebZmNFP3OsVuXBNUawN/bp3dEBFZQwHdSI/Gi15jgkom2jIht+0DEd/xEDmwitudi
EFEDy0TVY6Wxg+UQMT0whnVGd2dY5ygUVOWzihAvtnR1qoaRO3sLdWzNpi2sfH+PPUxxINyZntg8
ru0X+rJx6qLOo0+5oR/bZY52Y0lyWOPWp9dmfnIe4rUT7iYevNo0Dz3UEAvhacm9xAC3E+H3Io57
OdMjPaPIWVOV7jL8CnCmm9gQbw6bWxalW5Ej++jBmMtPIbvXqaCasSBis4abwagAerTnU0Pvy9rD
55OKcRWrKSvdTjF0u6DLg55StdD1qCGhMH2HxCzjjM93KyU35oFoWGQthQq9Sgdf/2DFFJhurWrq
nDNLYWotjqL7v348CWNiYpaCjSayVQt/Z2ZId03swhph/sdBMhsOBwdeHknW9FY5urS1qVn7wkjY
0nkeP2mDd3Gh1kwic2MfEMsVaFnQCaJp6dI04HwCopZ4n49G0yWFxteRbmyCP1HZcNZzlgAwvRcs
8ToCOeNs1degy+ym+UVaF8BxmUNcdYfhZppJf8sGPj9T2DgSkSuq+6BK43zCfba2N8wYr+0VGXnT
LwjB3s038caMefWSecIkXjVlX9+11hZc+tx3rSuynV4kIFYqKJs19Gd61vj/EIEj5QY4AzRF2R6i
Z0zHjFIuSTNh32V/eChLGTdGBzCheY7kDxQFPcdxj9GUULO9aUAWyP62jJzeAzap+F0LuUz0LmI3
JHsQ5B7Ps3PRW5QqBh8XodtC4e3KM7osE1yAOjPA1mL6bLGzb0zts/ipSInNKlHtGc0ADzq543R0
N27xSVeEBms4Mtk1rzHUdtDlm7b1EY8dqnjW4BHXYQ6QxQAIjIFbv71mFAIhyOWxSH8bxHHbp7bG
OoHCFFf2+sgtgwVtxZY/xiGJJrv/6DV074CqBvzMWrup6HuH26fmbbWhnnF3EaseCGcrH0zA4Kan
Rnat/Abiz8VSIiY0jw0uUGgp1lLj7UTa6zAcmn051lr90XQXc/zsb2Eyeb/PTULIjKJ6SvGUfzf2
kS4ZQyoo9IaTFRr8cgTvtOJXoKFJkX7yRYMgAEYtZAE7XQayXQgrl8jeL9YaSMXD2lZNTmr5bXCJ
ZQvA0TQWJYovIjORLryBKYnHBAblP35RmJ06LsGh1zY3SM0fq3bXyh6ogmFcEpVpefamfFcw1Buq
xhvbhmyapryCs9RJkpCWDVJQWA6k00zzO43VED/MVLC1JCm9QqzbL9hHKdhJecUHo1wwCcGGN/AX
T3qRzB5BWrQfZyHaiw6NO4k2VQWiMeManECVs7ZqI2qAOWwf9GgfaC+zg/DVnhGyD+rYMiZGFQIE
bWBtlM/MseiNjPFDjL2Oh/LKaKNESmG130kGtGgI5ryJr9gok2V+SUSusWVJQbF6Ez8bWbkevtwT
WVPbsdUZB3RabmLa5fmslh0ytbY5ut4eU1ZpoaEAfNErfds4bH4g6eRFB5PwWhsu6JQeK9ebrS20
dL8t2L3aqQPu7zS2V2nbIzDQVsfZfDqGKSxvtj0bJi6/c16BMqvJw1bKtNGH1VK28me4iM7el4i6
gHfpSL3lwwgxO+zCkMhc+xcv2n1u3ZpBI3B+NTkb0tcPHVndOC5jmwFulhm1aK1ErY1aAN8GGs/f
/Trruo8snnO0vpn6PXvFbi4fN7MapngHdtgspPcnQRPwdTMytBnHU8ho47AnLsumlJfwY7qx5VR6
aD0IqdLSvEGfPXkuY4x2HpnrVx5+mu9PdCboFqZO66TMvaOmWyQoz7eNkIU7c6mOVHFXKb0DOV1U
ONrk4UXsYJ+7a1HySQ5vuocDQq5CQmX5qq8eXyV0993C6wGidiaxXi4Utm7bSXnr49C20Piz2jqR
L9iy87S0xEodlWXS2unRnVQwzZrs/KeQcfXpXzV093lHN9Cw48J0ajtTdSlbA9IFNPUxwQNMiwEc
ruOTo187n+yRrPEBQS/rYOqCMRJN/JW+zKVMOhaQbJeUJl5BPChFaoSZ8vBi4YD3xCFeSwpNVhSa
ffr+cT7fUZvHcBH/+hVGyZFhlp72WjHX0tM7PWI/SIUUcbgJgeJ9tve2wjJgI4lbGXGw6lqjCA8I
mUw3oJ0uw+3SpVrH1xnXkTiSkRGx/y35ssqFth3qOQ/WhB7LYg2K8mWY+R9dFqYWaMoT0qFlml5q
Lfi5rdFrhbZl96kZnNM9z7run9zSEfaqXMwVoHsLrU9DG+akDUD+mSXonyB9nbGzRklrSI5I2AYu
riI0lHIeRESu+LpqwS8DGm2GLDwk1juWhTO6D2/+MWVxt53ruU62YZ8G7C4wcb9pU46d7ema6viE
VZZ/rN5nXq8jlp+cSeOt2O8wx83UFWAJvTlhMZpOAXN3uBKbdT+x3YgukvuAZwhh5qjPftFR71Pm
1yEA1vP5Xj0gzoH/yu+YkdwaElW7GPfIuFC1bG/P3QewBIwk1toIlUN+G/aJ+/yBHJJg1orMwzzU
FDB0kmmAVyMisDlLA7jnDlFOib1cWESTYgE5gpFOem8r0/irA9Y538LawmaND/XQsQmbqRGwIxtD
BUdPiC5cdnbz0kLIUtS3iZi1nIxmNcIy3Ne5hkHFAbVMSD+B312n7N/qEm/DyxdQCZKcRhFyABeS
Rk2AMDAU2LB+g6ZxWxJMnWC5xiIFQSqeFtxs18Ye+3+CbbFxMjEUryUgH1wP+hz9GIIDko0Od1R9
dkdo45/WRBEYBV7OVbrCao9nV2f37Or/7lAVdc/6g+DSxNyz+PIBfIId8U7RkJDji3nAIKu6v3aK
XBJRCCsBgvvwwz7xl7eYCDq1QNA9chlrJGBVqfRcg5F7mf2zsjpPNTU/bgfJEqDZavKt/fGc+qM1
OmsIhPDB0qyg7xkhhpw3lOQMguQg6NAKMhZDAavfC5FOjDoxVjJcNvHkWZG8mMaiIG5je8d9AxPs
lZL/aYK+yyzS2uZKQSRZsOcrUc5YUzWQtECU99YFiQAD9X5JqGFapKyb6+VXow0wazxTXJFRp+jO
0qd5Fhoz+Ky8Hze1RDtSJ2BX0ut6e73qJWanbDY/9Dax3ezfjR10JSeMTk/VsitT28dC/GF/45VA
bYcs7g0n8ZAjJc7Y/VQlu31Yo9SqoacjFPFBBretoVPHdxbCmNi9T/J+zibTPUGH8dYRdxjk5U2G
NH39nkjFE65ji2Rzj1mCtebvnTs1ucNgUniuxzTOC/da/7erlljOfRtz+KXw+PBMpVemkvuZ1Pmo
ebIqyws8XeQ3QulmyLwBFrT+UnBBzgEMnyE/ofOgH86Gr/BvlcpxplysiF/y2/NKBiTnfKZZo3qO
DgLWJZcArxWvVmwhYXxNhGZ+LKi0uQoud/wHu9LN8gosIzkouZQU81KtqTKN2dTAEv0Ccvm6ubR5
+6DYh5Gsk/ib/Cr7M/Wwwq58pHG5SSYHq9DgGMzfSsU5CeBM9qx7WNrlwr2fK/jXGhqehCRqaE/l
aPJgdVUoncanygx/2U4vpdz/0vhx0pRgU38skFvOuyNdMGhcZM2zFsjGIxahrJF657+wgFLscBq+
y4cGE+M5UTzo/eMxjrrgSQ0iK4F+KZChM+la5hHDGU9jjjuuGCkYKeyPzQjRbmZEsHZ1GtHdCnCg
fBZjPS5uH4bAPb8opqeFl2ioEYn3PkUp/+eH1T57sxwDufUWW6CODpR6cKugvROHnR/IjxQFMMiu
/L1s1phccRNc4cg5Rwtn/wdBz92yiiTVHOgi7ovsPQNu18kzxcbsGqEiLNpVQLUH2/jen+hadkBR
xZVO994lldW67SzXvwTTXZsk24kGPoUZCAfixPE0I4ktt9ZWhVcr7cOfmJYWkeYTJ99DzMvWdRwt
sxenhVqpiIuoyDIV8rw9OgVfH9LSszjuGfnYQ2k7PLsABj1NwY2TMSPBgzy1ejF4jiAmiFLnH/fY
66jpf7C0uWNv+rINjuH8mmrxtNHLZxvxzJ5AVxuV4JE7xCNPwnUUbXw3dw0G1JyRuEdtlx3D5T8m
w5yeTNA9tTYm3N9i/Pjr/YYmj/voi16oePobokpLJREDYeMPOKe6AA6C3O+Ql5T5blfOAAtzNn2f
z4oT53wGOz45SYlN5TieUeLkDwcxmnOfGtGMNAh06ozWO205BMTlwzxczN029rBn3jsF4sqa8PUJ
LoCvCnTM5fnrOsTa/WbSQt7uBmYZSZQdHZLQ9W7njfJccAeOqk//0LaHnLDk4GtGQdcCFnFNfg8y
qlOkHFTvMXY/OPsPnJ7XtdPh9ID96f/jd8nkaDP1wAXM6F13zWjQgnDHKRkMmPIPm7s/WTfwkxDn
DZ6xwuL7J+jjLkfSKlmo2qap+x53rpJ8QzK5S/8cAlRTfZAIxX5vjo+VR/HlgqzC8HfrX81l7gqy
sssgl2Q7U+nzxLCE9njY/IIU/BV6x7R0YBV7lnwikuKsbTgvxEZgWJXh5MkaRJSvczl2vYBwdjXw
Au5AIBde1OSTEndUOLiGaPPFxbdtWjl69vIsQqV2JaiR85q0mCeaFpe7A/vjx68UCfQCyS/AuNkT
Q6Bvsyc37zk+gKxrLAHFP/i+ZKExnmlu0DhiPIBbnqdXJ6008Dz2uV1aj1fPfYWdLEwdUouq86ba
pdTiSroA6Nty7NvFWqhJ/giV4oh30Ba9/KruHWME9nU3CHNwo0IWMLgFsOxo+55g7uciyr6iW1Zm
Q/GcYFi4QJNR5CGMOOzMzzzYGc9hdLBbT3C8Efz4GcQ+L9zn8h892U7Fqp2OrbRiPu09BlGhN2fu
cKXUVAfEJtTGF5DifcowMLk0OdFiO9AgLzC0zgQr7hOCDmrqxgif9swvcCv6msTOgPr247k/vNS9
+nXBApWPnVMHf93/qaOxDG/qRFD80K7M+Ad7si8NGrkrzHWyTRu8qv1PXXxYsl8TdCraDFdb/4JX
GW1ueMRYmN0ue8mjZVNQsXlE29qLNIy+a4BKDIoSEV/ZqM+DGcsj3f2t5pDrtmW3UgcNfRbypZRG
5iH9k/kxKADWVWJxBfaPGE+kgTO+X3IGpRrErxX+oibmDPcJOzTAIGwIEtD90rJQRR4WHlrmom6X
PuBnm5OJIO0PWkuxZAR92Em8POfkZw41HG7+8BFPAKKHJGE3zmhxlH7FfOm0IDcpo6amYmf966F4
H+IxQGkIotm55Z3B62oRc8/udYdLwkj7n8iVrQwmOz9HVMkOWfnE22afFs2hYXxCvI1+7nSe9Nql
zhfHvV1pF5P7BBBGFIoS531gzSa1ryUORLkqlu0OaPQwepS+bIrMduah6214ikK5NmOJefXvGkX1
2URvtloIknFzgUhXRK6y9IoAO0ElTiHvm2kz7p73GjpzQ8Q05Ia+qjOPabOdNihcAvIn4o7LBBUs
yAkYxBAeRt0TApVQhkzPtWRlQmZq/j3cdZCKFDeDCoerX72KmnhPZTbasRNqcc4700V7t/UjBC+x
biWVrdCGfMEeNp3PYf7wn6SfQE9JzsCXPX9yKu6LLbs/3UZwdEiDj68o68TKenSfzQx3HkNxSyC+
GUsc91r/x21knLC0d4ew+gTqfGcP/IEWoCVIgrCKzpJJTMkFwgS/uT1rHjNF6Qh1yDSh5WTG4ntH
AAo68PjTrRL2xq7wejbtyyljqFlTlIjwD7VkhH39IdNfYNllOF0rHl3I65o/XCG99Wjr4nciJsCc
FKdwMBIRhbm+2VkuvdBNgnwdLsQd3n/FmPknfl1HyNEkLvgy/0Q/yE/EFIBxvVTEA6DEd8bUkoZr
wfuXKVRQ5MoK9oSgAw6Tg3dYHEkWdSUkzHqgQhClwCOAeOFL6M45ZKv4/ye5zMMmH1d+AhSY9nrF
qJNWr+86xSS3N4OKSKzaaySjFB3jlgBz8MelLb5UXezL2E4uxV/BFCRXnXPZxYNw66JmHU/jvGcJ
2pzf4ZFkjaV6EuEskclmVRcgFnXqYPwsaFSorS4sl0j3Ea2YxT58UHGGo76yJpjreShXiH6JkGoS
rbr4YCGAC4eCpfCjaD+huSpbILAu0CA1asbXg5/fWXDturQ=
`pragma protect end_protected

