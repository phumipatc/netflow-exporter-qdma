`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TJGJcVGoqM9qzXnXITcmmQupPFf/Rmy5cv2S0AAWWTjloSqezTQQBsVtKhOlMAh/ip+ub5D08aWv
+0QwwoOrKn84BsybnciQ2hARNv+1di1NROKMpz8N3DL0CVVH6mXoybooDHwTUZeawDPzBYHKtF1v
qlPBDkTiCZ5g3ujFp0jCQFalfxQATGemDUiAh6mx06/6nWa3LtZ3MznyiT0K37xxFCNHdeLZa6Z0
W8P+fQ+a+1ujyMR/+QoYrjhnDLgnflsu7/2vtb9Xa7c75q4A9Oy7FgLxocfd/S3qycs2mSWAWR2k
ED9vJkOhe+Ff0hCnd4NwqT8egNsXeUA+yj21EA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
cVDozfFRr5EzuUdOZ7IsU7U8PO5gQ/oiylxytc+BVJyCi2rr8bbR8L035UlRmdwGhf45UO4/qlK4
umiK8evVakdbQrPQKKfxFJlpLyKonh773nf67DTbSKbAg/GpZYNq45rsFG9xNRpMTeAdzyzjYcxD
7rqhWKsVdwHIwFDbSev4z2HFfM7MK+06A8vBs0ytceB4sMOeQ5Y/uyIQT4DRyMQKVyoANkjxNlCS
beqPQILB8cY225qTxcUlryNNOw/mWL8X/zpz/ElJdgZQHda+Q7dHbIqeeyUhOwuu3Hd1S+8S+IQk
nqATOy09cenMiDRYWaedpjUqhPN3n5a5bafaAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
pwkoHnh7hVr4lYpWAdJyeZPBy9KpnOpe9LJGYfjQ/RFUE8r1al3JvWdOyw6BXFjM63T2VaGnxFig
GPSBYp1c7Q==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bTkimdYWtt4zMu+7Q1702prDhEns5RFpVEbgN8sAxyreU72pjrbgR+TgLzSuXcWATBzOBbWbWagB
RgYsACVBLpym9fK6klPpIjYLLmj9O/Qbvl/MCGDperWOOZP4NBZNOGgOgWCGlDo934VMVVH++Fod
HU3pS3oeHvghhGwSz3+bSob3XoYZYj+7TksX4zXVLORK/LbTiDZA5p3UNIHJkf3aHKk3V9QI8R+S
QU2IQYhFRyYvwctvwW+2xqeHNghXdTUmZq5/FZwwRJy+UcfF7U9bhKq5gpfm0I0ElOBGDWC58POv
kuJPPTUgt5BtEM+UW7bvVPpWaiefH6qyS4LPPQ==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nAIqG1vX8sPpHToHcBsuYmJJlGU9OeVsL243gIwIpzjo98KKD6NG90lQ7N0kFjUIfq78IYtMSM9y
yI92WZZkC6jBxj7YatxAcJYi5dMbyeO13jne4HEektRZo4YVVARvihKHxEF7Jcos8DruSDjnGxlt
hA/9abxJVgWW/hCanFQ2RoqNuEHFVBha8lgRhKB6cwcIxHQxGgt7K23lxq7iEoDBq8N6d04v8qt/
yvo2KAFctJB9vTwF8C3zJ/QSrCFjxTgrUTKa9yU/O2KfPem8BVYCMQN7e+sFV2bwUXGMmhnHAB+Y
nTDr+cy8MW+0KLw5TTwUhkkOyd/hBH398QSgRA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jOZi76GIXIb2ae1zZCKYSIJP01q5isHNNEmij5gYZPUgX6IW68u+M2tYtzZGQgTqZmaU6dZ6iyOd
61yt3HgGKIOR68b649f9IA+FE2T9q2mqCOnj3uHMnFe/SD3XuwmGojmDDhz4tPDHCFpVeZ1vLFjH
Rgx8HcRznyCaKt+VT7g=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
UlvXFUnGvJuzWQbiBvm+PZLvu7N0wpQz9SOxO63CACYsL42jacrhhZJsXyQCQ48VT2yjKFo1cODS
2uvtqM62GdlJIia7hOm81zfNEIsuZmZBX7lPp5P0F/yCKEZyNBR4pVDLo2rAvxbQAnTkuJ3MBYBE
BxIRejlV0793ZyvgrfyiC8WbO3lhdiEt19ArNpC0zMw/Ff/NUlLBpnIZjv2O+u2V2AD1wVGJgtF8
NpMOI/k0nFAUJMrvVYRRsHqh4LGdBys18kGU6u3DZjOwmKQYd82XBy7QqjAbkMWoIzC8ruZcWjZ6
EEfWPx5lhy1on1ox0tTSv64LwID6JkVM7VrZ1g==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
t4DaxFplGWEtwfJOypJE5nTfltKqR3Nqf+gYuhjEKbNGfbvyEmtf9ckiIImQP8KxYJxDdzDacQsp
d9OJsOUNL38kKDTlcdgtkmo0q7KC6GqkdkkUZwpDoPBjB1v+ZI1H37gV/XGM7fFuSMzoZH2TTPIK
+UihVxe1035gSJ5+v8fm6j6pTpbBi8XRxFz8O8ftFDUqGOeZVo+2I0txGT52/XNoTZBMyZ750D33
Wry84cW++zqJcEWiLM894pRJW2xKhQOoAFbh7+FcU5E7bvrgjWd98qNQM4F7tWcNxMySCUBR/1D9
E+gVNZHC5gHP7NAjxLxqZ8d0EactRi1s3pLpRg==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SQTapqCeCQUmdXyZqGMlQ14nxyEmJkERK/vqAgS9ahck3JTut+gFqWQe2z1scriKTErlVQcm84Ws
FJTc35zSZqIrfQ8WVJO22fi6+6SRye9m1urmxUCUZUvB2EIxBlljzGGKrsZ3DwEopk0puQbYIHXG
9dmSpP0ofChNcRu4bRc=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kZL010dI0P1alftVxSOEBGzSyuIVbjGu9n9J5jTmWnPwa1c9AirdQAI/Vrc4AgX4nFL2sjU50k+2
kMhtIcgXRSmP270we8DUdVvkwEobygQ+N1d9/+9+F1NklrFddHGWdcfngpQSmAxl9BsLuouryF7F
Xw+dF6PSzct08Ev9UCE9Od9BF0XO3nz9EPaNvs9hw4+auf5lMERhog8e7uG27Do0Q7FLskhfXli2
9y1twYGKJE9wfHdH91Nw2ATphSpYdAWMsh0l3PnbzX0XoL4xv+px/Da6aaxJ15TA6GJW4BgJ400k
FyiEDiQ4WcC+Io1kAVyqTt7uzHPfH35nV/HegA==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36800)
`pragma protect data_block
8kj6QeffR59Qcy2gQFOZ1MOKnbveARGPtDknRVpPb0TcIV5PoBQcwhwWvp6a+yXvgiqGZ9bpT3RC
7dTpt0apoiNte/qM7LQFszTuV6PRy1rkcvmzg+TOYm0+N0OCziqFEpOL5aEynOyWD/0Ld5HVFije
o3kgO7WN6lKMkUAuAMQ0bxZVR8VxZBo1PcwqdtUCLVSV0kOxTWLizvHkl7nurASLSsGq++Mya4Qz
OTC3qj3FXA8jX47KNas6LqDD8AxLNFxVXeq1eO1yldOhr6D2TYFMzolUcUQPCqSWSfhOhK96jAdv
sl6J3W8H8WTFE4CPyZCj6hZwiQ6NHHvmdeDK7gW8tvWuyd6J8odgu0r+gAf77T6GQBc3zXUxEhD3
SgPzXS3lt22IMavzC87JGvaqf5BSQ2XE7k9nlySvaqPM/NjuMRxp4LOD19Gukz1nji1QLraek+v4
hfehI3K6nrzOJAVcjXLtR2SjjMHZ1xSdpzQtsRVauXBg1lD3rNwck4JqpR34hu2JIBJwUVQgqxQ1
ogVMRedo+tTX3S+DeRtYRVUrNHddBp9Rv0ciQUaiX/xgfeONHD2JCxkNBAnTn9iLMFqcL7kaIH8w
b5hwBtMoEXFe9mKHVnjOHIiO+oUC/bvbQDDtZx1gm0RvLwz11GvichgW0kFxIbhTwWNTs/pYeFCv
Mt3Wr7IWYN6EqQCd6x3695Rk1K8o8zgGLkX8fgbe15Dplvi1GWFTivazbWtsSD2P1IfeKi/xzeQl
BiNQGlWOkeJRa2HEjGEczmX/1EQ/9G6vcd7W261RnzEx8b1LJ9nC5P2PizUrpB+KCGlUjU3qT2Kl
r17Tfr3Wwv7EhYtLvP4RZgQwg+BtvFP5I8untUHeSEHRyddQXphghPwIkImG/CaYo/st3zSsPepI
LD4ZtWA62ENfVoDw2V04gMS3qKqYU78GELyueEtsRKj4gpvflJYFZZ+UAll10pMPiSRs5ecn4Alh
Jk1VcgA99+QQQLrcj80I6VVYWaz8OzHo1bM+6YvKg04Ijc9Xx6ZsMO3ED/yTNv86CJnpnaeHp9Yg
ZVKw85R8Rsa7DYe/d7MBA+ecvbhigzrViabxzTaShLO9+WX/b3MJa4xFCPjxtBU6fRXnLk1KjZtr
t5GbDBsdTj4GVsq+8Fx1ijsBGQ6+oz7op7gzC/z2+AQ6OGIzCcL5A//V7EpaptvXA85r38cYIf+3
XfldeG1RFzQ/LgPgzH8gSjLRUg9pquB5cL3dqkjMVekPZi/mCRZpTUfzONnGVBgv5AIm5jAzLUTx
yGRD2pGhVdNYcge4hUxlet5Zw3lrGfT8OzBfEJy2OBkRurtDkj8bhAfn4Yw6DxuVkj/W3kpNnKpu
/W5oEuRaFrQlz9IefI1mnMZ2tfH/VBqyK3RRV7hHGq1nuW2Fa8jziWRI0paqQk3iFDaELZQeoakr
L2ZTg3gm7qUmzS9h/ydaqGKKIwCG3FUx/4V1WMNSBIaQwjTtUhizCVyRg2jc0YkJ42S/ypW75PBK
4073YzDp4+i7erY0gisLMyw4j92Qeet81mYf1SUeDE58s4UIJrirIEVQtN3F19upUdYlnFsIy8K2
Qgla8o4EFBfrW3Mv9ecpkefKSbrM/gypNL3SmjPFn4TsqV5R1nJonjnIRtAQa5iU2hz5rKAd9MGo
f9B6ulVjlpHWKOS5P2JrOFixeTtS35q9uk5rBa9VDu0U5yqtAHpkF8N+3txK2p9qyu3HnAIqjvgT
3U3djp32tkevOM3vpHtWUh+p93nzOWh4WpuYSGniT3JzqkNnlM47ComRYiRG9qX0kZM8JolLlCnI
FPJwdq4fm3HxnIjdtXif5UUFroQwKYRVrj2grRYvojpPlp59pNnR3gLFF2Q04aCATPIiQ9smaCES
T/O6TFDnY4vVuXHgeBmyuWC4KOYTX7ANQwlqcv7vAvKyagSMUjS0JK/LVUQQDs69i6mDb9s8S3w/
O7eheqFxeuVzHkp0e5wl20Ltj1sXruWNiVRC47o/12GGA301rcuZ7vKddl9fy6zYg3/PzczL39zI
lovgYFOWaHvi4tSNvK+rjSIQGvYQdbXmOMDuufd2lvxsAnRjN/3UFT4Ptp3OAXn9OKwWZ6y8BL8s
d6RHtBvxzXfNGlZpNKtou9c0bnRXM973DUmoOsqgPX2kknjHOtB1YPG1NUMGOy6GTi6mO5HaLhh5
9JgbxeHDc/aPi7iBbDmUeHvNxbTDZZF4A220etT3cpwH8/j9zMHbVkSWsMs5uagApXdyCLIgG+qH
p6GIFIXKp5SRx1AqQCU0BhOSxSV1ODzEv2XhEonSlzjk9RNKtsuLq/5zYMgFHPnMO3PrEKhCjBx7
PHyiiVQPJ8bDp2CloGVwIq//uxn0nhRxCWVRweuEpK455u6mWZCn0/yjmXTX62rqx21+CwJHwjSx
fMuOSytlemKy9kJcoCIrdWxIZ68sr0y9/QKjegfmz4UOSanKxC6uqnLSJorRaGg1TGyG7mXqce2A
3wVo9O0FdBljCXbl0Ofl9tOug1nAOCvqDrafWZ1qHQE69LIF0lb2qWZQjLTXQ+8NZHXF2YvRLsW2
0zt8xp4gquh3jXQ5ctJP3GzT2TuRbGj7v+j1xmbbiQ3FwFy6279WQ43vqOjqaD0Att19/kR7+c1C
uskwwgdCzg0B4k5COueg0BdIODRsnrISeoxSl5BSBLNaj5On+JxbigRKLLqRv5c3zFDa90pdT6t+
X3aFfMaCc8j4gb5VbPhjw09/u2HG5Uibb5VBNb6p4/HEMZoV/WDi5Uy+1Dn8VooPzUXK25Ojp0GP
4D99SdfLYfeT/K/w4ZhJggz5um82nHudG/++K9zVY4VtxVebDwW7FhWX6JVIt560gtAHgamHdA+R
C2WGmalC1hU2Hb2GyDc7HJ0ccU6XcSDdx3GqtBGbXEh/cgr0BnRRJI138h22Mm80IohJIUc1S4pE
dH1UBg0PjYO+lP7oGvV5rF7Gq2RRVPPcQNF/blCMr2M4HHIvHHC+442XZkhosAFRL2On50OMiVSw
dAgCgKpmtcvvC+urWamh1OzN8EeQeG+P+Ygsmday/yxubb0nVxHKHk3QAJ8KUJN56WD5d/iGpFGE
mk21QRcDDffb4GOT6NE76v3ddKTNwKiMQ4ruPsjtKHgECCMmHtk38GR9B5id+WUvU9gTdFNQCq72
gOB3b79cwtdAjWRIQ+tFGOmF7HdW/DgPxEmFmEn2WkLy2BqqyK5ACJwAmS8OnCzczj4dVonczoHr
nd/aF8Tr2lhK1ZAZ/k3ULWHsACufcIguWeItFXIK8wSOqY9jQoxIughFaoxvwBpllhjlK9q+uShk
eEdaveDYbSYf/tWZghmpyWaIkAz64kPVu2osbrymX4yGxN6sSPo2b40YrEtVv4RrrElKmeb35j+Z
MW72Lw84zmMxedU37xo4VzLR/mqj14ET8fyKB2JjJz1/hUbZfBdk/VQSa0wF1yfZxGIdL3krhKoo
Ewv+IWUcODpX/RIwsYsMLQv3s2I3eGM1jZ/5M4InSKry/iUhWGlwp+EK2TsIcsCzfTMFF5lh1vJJ
zQEKIKRTbSo4zSMAENGTIS6zP7Ujboe2Un6VhHwyn+qVKX/Ds4PNrRpBhbVJXm6KkCdtyTzISmId
nuwh1Q5wRHZuoixBsHyTaBWZ2I///YVWk8k+yRFUMkq7/2v7X/03sJMQdIQzZ4kMdjdnyCpvUfVh
PI4RWu/BKCYw6gY1xs1Puxy/+pcE0fbAdRKwkA733T+l7qWdgy/RLPHDv028sLs1JlEJF8li3D+m
5YwL9YBZDRtpygFm+qQQn9aN2T8GC3ufQJX9iEN3CiMxxOPFRgtH6nmjHPiFAXj+XGcVOMDQWcaG
M78hBZG85DE95kUPBmMyx4RfZ2RkmRzipRPHT1jOpA2YosKSCJMz48TcaAbZiZlA2VnoEyJU5Kks
GbhGZ0d3+A2uvewKWYGe4jpnt0KZI+xjiDiBjYeGvKNDZByIFO11WqtS/6V4krdYayfpMIqGiXvM
yUEP7sR74W7CCfqjgW0p4an7GrHUvMVqDG+BPf9Y9fVa7fP+pJDMnmSnJx8Q4zMO92PWmK58znNN
dOS/uVYs400ar8bshQ6CwSuERDg2+QO9Kr/io82x3mJA8kiPIrZpr4GlD4d/KItfJ5ry/LcOx+2X
oMi5uRPEZhE98HJfGOsVtZmSiAkfVAlPaZsaIXnVizD5+RRY0NOAyOHRedjfOm0dbFVs8QwWMMwd
YVFn5iRnmsVmy6MH54MkXtMgJJcEw0ufjR3gyyESYR3QGUlP7zhm/UL1MFO0UvF4SlapWHUo4dHI
UQrVH3kqa0RMCQZgTu6YA6DmDFze+6bJ7+e2Ktvbgw4r/X5M1e6yvU7K4G+LA4vYZGmyr/u45XJW
rFowMPwznADGecUAmnnXicHVgOWYfN9wgEb1aV790BRzdExOr3/dKn4QVPlvHOKTTuDmf8Z/uLll
PXdMCqbgTCIArCj1vksSOfnXWkhuk/PVieJADblBC3vkhjcopbMWr6cs+sA5q3evVV8AgYpxIPtR
QvQGCdwP2kUBQAyvYhVPd2CzVek1TwdSOG/WcmXSYAFmY5IvywhwmqvWhqfH2RRLukS4GTIyzWDX
alJf8FF3K7ahWPQpH//Wg7q05xYY7icMqi+MjXWfH/upoPA0O9d764SZ3MS0nB9fJ71pMygdXxi1
KaE942N6x15sIW26jJ9+JCNl9fwNT1Ig5gWTO4cvESF6gsV1T93R9S4ZTMkQtQQ5RGl+YeUF4Urn
JgskYzkFPQgXLUJ5uaoMWLSFtZYJgpwfWBWUsv33FdkOfI+nlGqDLtM3zgJZ+QWU5t1Fl/Cfho0T
WdrTfWbsRLFtYGBqAv4N/riKqgpGN2zNx4mQIH2BRLq9sU5QgpDRRFUlAaOdMF78k7bI9yCk6VPW
9QHsFuoFJ4400uIvNIZBBK8WFxQ4A7i2JqlOB4/lhtQpReiVeFjsGIvjgJcW9XG0xeMU3sCFuAme
qKYmug1YrNgscXRGZgtiBndNcpx+RMmoGOqSSCsBgoOPEfwZ23bF/9GxgEkDR7REP2t0VujJov4T
vDqQ4DEKwtGPWIL6LR5MwjAXe7K8RAU0tPqWFifhwCzYXoe2xRkIn7z8ehXnUEO0FW6ztvKt5ikn
E7MX8yPjgoVEAfzyG6L4NakwIEczHYpHY0uiLGaThppDbTbaWaQUTyl3TCPwH7/OET7EHp5UrbnA
aTk8YrWQ9sLp51KD+IW6r3UE9zUVsU4MJC7gyBAwaY7jConEKlHnCZgaBCHcfzCymas4CHv7rh0o
m3YFRLr4Rx3paBNPsgiqYbPCb3usOGv1aSt9dfh5tLa6BpIg2mHczoAWusnqsqQ/ME7c7NIgjtTN
/95aMt7t3e9unnyJsJieE8yBYx61qTj/zfyKFBnEP3yzTMexqI/cFy3n6l2j5cCX2X9MoeThcWbb
MDEe7tdaRiXuOtA4wGTfnWsS64tGIAaowbuqNhKnBkkh8ZR/VMq6adzv5tuuf6TLY6Ph66Yj9EA3
yzFFV4QXHar5+3/iKv2Um9TiUVTC8p3pUlBwIPVFCv9OQ6Gn0KzItWxYKISQrZTWI0D+GOHxyz6J
69PhN65BRdOd7AL8wM60kT3Oa5n1tM6YhURIkKlRnmuYLrviUuMo8UViPvalhVnB312mtzg77oN6
JK0keHStzrLf/9Ry8yfNS6vwfovUoeW+zC+FroMe8DWRvpMhafGgvXd+6xntQ4GlWjCe6aklGuS9
VrUSoSa40w/uiW+c6YVLyoIB4kiMd/jrEtsFSO5kF6YlBxcOjtosLfQWJNgWonpE95qK4XwM6ppJ
hgqT23n+UJxg+lpXgDl/qZrAWIBT+h4W3HOegEkngl7CD6flSX2JMKDf60J9oClDEg+aai5TD74L
6is6bOVEpYkS+zBNNwyP5oWDKGVtMa4W4+6ckjl4lcbHfdtnXDerO4GzZ7OTuyJ/1HQDh+GrYpQt
wpRvb/ofJE/5+ZDVkDVyNiWaq706lhOcIMbFDzbinQxcSx2z/hgpIUHQ5ezz2lwou6ttjaD0rIa/
QCOen+8DGyV5Mwun/+Z1FmoUlUDfYkgJNb8NmpYyUhZfkuY8WVuU2KgWGP3Z6usM+JZj+kRQjYbb
IAYQkuxZ06WwU1YlSskFcdSop1kx3iRpndLPkN5HwhbSj+d3o5fuDFGAMSWkeiyBJ1/DNGfhQK5o
O6gdlsL1mvGSvEL2OYu2Zzv+5lOszEshc4SeIrSKgyJPYMOtwo+o4YSLY1DqbSykXkWIPwCOx8Tl
u1KFiXJySNaPzaHEvkQ7SbDcg3/Do46RpJtAXaUnDshZ7e81Y1KprqriFeaEuMWb1IucZIaIFY7j
xWhjoF5EKtqTDEh5NDPJLavg33Zo1A85VkTup4L/HwWyqhin/xyfrUwMFvsDjXm2/pHDv/Nx/lDs
p+2+D0hcGrYWP+/JdLV6R5sNBEZQiwQxQB5K3BPuJ6ezgZvaBDKFOwlbKk0bkN+06khfKlKECM+/
VvXoiVJGMc5UgoPWKDF68zDLySwecaDqt9ZJyBKYknLWGJrguov4EBmErRG8YnGWHOwWGHiozqVa
s9hlVD9ltSfmlBDnil9srToXuNyMzvEoGBdfNlLxg2JkgzP6EJMDuHIBQuGzEey16UBQj5AmP3Dt
Q+qfZZOA1+URo7dp1dCozphhjrtCoKSLZgQQNgLqEZ88UoQj0SMAzQbFXePxy/kev6YQgmHXXXuW
bi6CcK5ovTxZlv65n3Vw1KLbAdfo3LeoNe6oHlwpmZnlDXqQT3UBi4iubOGMG9sUGHLkSkgm7XUM
eO2Bs/N80Ey90PZsQe1qlgnW30SNhhKIUTYO+8n68gancp1Fxn37Z4SNdpDKcPs8aYBUDyX8kUta
iTUkmMgo4jC/gUyBUwgV7UlW4Z+CcqV78e0cJltBWi64RjctIO+17LssHVj2ysMi2Z/H8DkYJa25
OYxowEzLmF0DUJes+jUSgAsWv4cISUrJeapUgPEkOLzkEyMMdgC7S5PwAcXzA5uEL0uJ5OjkWKUJ
VW13TyY9VvRIc3XtWTTUxHplfONrupD+KzPOm15Vx0uozLeYX2X5rhLSl2gUaignbAfdV7BikvmJ
ZdkO055kK7DQPZFjTNCR5fAie3dhaZgNltIWgxuspHjq9sUX0Is4KzAFHpLnlMtuSpMxTeX0hyUG
vo6by2SjYbcllorbOIH8HXwBR/OxFPlYtv04zXysrlenGiwcrXAsJ+7sjpsn3PXOulqo98AWJKTb
7XRediagB35bHXMAIScYJU25kBW1W5tzaoWj01A8BGvk5SCnZevPSUgjxcEj2nrKyRf7C1k8nKFw
j2Fz3FeH0FcHdQJ+JvDRgSWFvcjzx3vKo2CjzZ5aV5gS0NTgryQaOEPdLxfvUyq5FO6eF+9Xe2pb
E8m1FmgEOaWDmL9BK0eFq7jpf7Q9dWw1gimG30qHVVn5oRIL2+9tTxSio8zt2zLmwcBcfNWZGfbj
2KRKk8Kjm2SeieEduTR6gcHM36YCMsaxCDmXRyqxtrO6ahpWk8oDWuLIveW1lmI0SfaEbJ5tFVrx
QO9oeUP1axYt9mbBTRf+b40gjROLC6JkKJ3ymoKZ0+UxeNN2+0vVXBUM/hYbW64n1gDUt/fYUgiV
81iYzcdVkm4FT6+5yh8loHCuR/fnJP30i1TwVG6yzYXk55mwpL2nSlgWJVZE2UD+Dm4jhts5Sjj2
SHtpiBE5L2a2pOhblzrngst5lsagGda8pz0aP1RfLjc5uRXjd9wBMfCDywy9KhqwhE9h9eGQ0NFP
mFAmtmkpY/jJfY+AEd3b6GIeuY5iSpDAkGTjfbNExeYjvFri4pH+Ei9wVtS4IUvxQsOOWQIoiCtj
M3r6vnPWz6aS4CuoYkQUEEqptMOzs5cBWI3Yvd90/6J2QYVEdDVT4SpT5oIdJw1ppoGEnZ5ZZS/H
PskP001dQkTUDcK1+MSfaOIUcQcy2CDSXv2AQDUscy+ddT6834TeIHiCXXSueAHbscHln+IhGb/6
wZB/ajuEZeOizvs+FSEQiJ+iYTDnerXqY1MkcyVA43WI0zohghagjwXxkr7yTpz0LulZ787/8ENg
tDWgN+0dePl78kntECnhw/2equ5gDgMd5YMb2M2miQAgpj8QDh7UUXJkBwNaA1rz9jc2lbLtoF1U
QA5srlkkL8xFc5bZ/B3yRGqvI9RYmys7F1QaGV5YvEl1hyeoIpZTA42f0bJ2/YbKCaoRhE5+b341
e2f/Mp/nkuDTxr5a+F4Dv2nWFE4ZOc5mXeyjtlZl7kSUVoI9iNambdALVv5CxkRjUZu2eSxDmTAp
1SdURDQYK9ISh/EYYM+Wf88fTuolcdFHhiH8l/a59cE6k64dPy7O0cPz3JellsVKwXs8m0X11al2
Oi3vUTZIVRH/HXzRB/JYn5GZyqiCcIfwT9tymc4hZJpFPHkTX5Dt/Aw+C0Aos7qUKn7JwV8BoIhh
M5Qz0vcc6OyV5btgK0Er9Vh0PXVpW0v+DTTS5HHsU5OTXCkuzAsx1nCKY7b0E4gfou5nzgfWG55t
bYSljEtI82Z4BFyTdB5k158KkXeUVH0BQwpVInRxDjZRJkk9wwZJVrfzKk22AalsumhgBkdHtP/R
LGgG9fv2gcJVBN2En588n68D2WY57OP6o08g4pYCsU/e48+EgZBzzXF110GDxZhkUWsp5CdDjPIz
hbu7kYxPdsU5QC3EJgxljLb/jyH9KBV8+Y50lHxw6YekIRoxKkLCOv2ywbpc9j0Hrd05I9/D8vH8
p+10XBbmmvDLu5PXrK5Ztamo8Loii9L2PljCQcuKUv56Q1f8MQwlHCzrULXWPUpRuXM09DivkFhd
f8fYNNyX+8a2tVal1cg7RwnFnqmvQfErGd65mntKpBxR0VBTYfrEF3n4eQy/5hyfC/UiP7nzM6fY
m54AsuqmbJsYDMMUs1JaNbuDLHvuK/rPG1BiZWic7zSetNzgHQLcdkY6onHd5tl3knhrHQsdh7oF
DpgS0oj8SA83I+HLedgJsfesfqWKtNS0N6k2d5ASSH1AJG4ecCVB6t/8WC76O3nJPCLOGqR6hFfj
uCMN6lmVvIYN2l/tphL49zyC9h3kqdTk5w7LLy4Dxkabxb9IQKd8Ovseql4P1+82Rh88RnAgGTF1
l+w8iJiEXkehMdkAiS2yx1uie5zJ+28Z23CbRa44PhArY9tm+A1QmR+5qXZAeAV1i7wUYshRNcw2
JRt33XSV2js/mzK49PiVop1rc5u/1Ka/JwPBI/f3a8+sWUVOlkTaEPoZ8rsyhIQttP92uAhzVKsW
DTPwva7Tj5edjbHKXe+UC7J4jXM3Fa+yPJh8j0p5iAgE6JM/ZHCZYFL/13ihNidwjaZ8y89gh5b1
5Ax521UST04h9w07hNLmsC74fnw7vPlUhOzLR8LKm3J+5uUsauyLpmAXOlhVbUWQ3YBsyw24IfhI
sgQK5BiwmrqxfqQGjN1imII2GQqEveZXiysWcM9DUMD8mavr55zdD2WZn9gzV95zYIvMXYx8mkAq
HKFMKLRUyUBkM35lS22l2mncjdoIqKoz9gGqpIk3SYeaCYuFpKzZ72y6DHP2vlEEW6R3HzKUnl0N
fotoYEjNSk/9NY/IOs5XJp9FzZdbCl2XfqRSGZX4LwBqmhc03zaJvSCqCbxsKHWbVx7Ux490ERS8
n7Dr6THmXdYj+0LHCb4bxEMPMxGXhJw/R/ZZgb4zicHJyeC5Oe1VVzj4/ekBXIaUGsnM8M3ABZwa
7ifdsZGh96ueW60jWZLbl5x2ZJ4H7JlonBbv8yRbYkXgteU8y+yCBG3HSTRyjHssoeRtqQUK0m6L
zakZejfVxqNgK4zgzHkmKt+6uHyJ1zhbOabJTf/aPTDgBMaMS9t+MFVKcBCwRqQU9WbMuu5JFLYg
7KB99kvLVg1WRurIGT81yCZcbjLhTmbkFVdwOIl8KdzyCgPf8Wv0O2BXZq3sm4mt7lBv36YaZfVa
POFTf7RDTaCRLmE7AuHEa/dQmtL2XFSs5Z3QBj4yAxDEYUEpeFRANVAuDPAsDSxH2HQCv0uqxJKE
goA6idBI7b/UTb+BueA9LdO7j7mL2PqEa2gWpcCK4mjIp3xqvszbSVvNnzyu0oNoYpIHnOc1ZKOs
UGAK8wiip7ncEZGqsN4+HPuvXzaHb/ev7qET1MZovpjnU5S6ii1SUpA/mxprsez7eYICVu8qRJ2O
1h0uUz6MgFHFDB6SN/pW57aESGOxwI/xP+lQqxmXI9F9jXoZWhhOsR6zoWfS0rV9oPRtBw9K2kXg
vjal/rwH6tdOvvEC0xXSaNqtm+whr1rByEJJIvHgilSxp042qLo8NEG5OCYcDrnphBvcTxRR0x7D
rBvHc9NsM+JSjhiNsIQ+hOWhvzdcRK6Y7ykrkuqEDK0hv7nYA5HF4RcVNN7jge0MAN1BUE4mUGZh
WKaW1Fv3eNfuA9/QP2EZuziUPc7hoFp+UgWzhBhiYws8ZhloXie0bhfvDstlKHPL9MfaIIaPq/6z
LchCooWA2O3dMXeM6j8bg4by8A8Y66A/FnMKQEjKHbUlC5YaJXZXtbvYTWuNeRVN2xIxDWMARg+r
Apdd5syaMtv5YKNKH2id+O9YGjs/gZwG7ls3GrARQheFBHJIy4CfNrgLu5BlOur2Z3+FZQgne3s4
Vc+lHskMPu9SAF6RRyR7EOdAnrsnRXIA+GSsHp0sh03y33N2cbZDuK89+BGgOvHDgonL6xonQnxb
A74PkQi3yxxNe7wQc+849j3RmLyc5ooh3RRLaW9ckdjKIkrAG44d2xrxG0jaDrHAtbzo9iUWj1qq
ExCujT412DpfcZAGoNgqWiYmpqn7CSDc4TelcWaIFhGWdQq4GWfJgCa/TM17UDvdvFkc9eX7dpkv
tHPvF5lMaiQqJHVoRay3faxti4UYG+PA7ttD5LpEN0WZW7pLG+72PuUS6IkOgJKV7RUGzs+n8WmU
jIJDd9cPT0t9v6c9iIvIAtlbz8FnOBS5ndD5VaW9xqcgL84MPslmM2Z47+xgVz9ohxPSBr6jPzdh
JkIE403z42/leNUrtrINDOPyVvkmKXklEVpJ1CMAF7zBXmfICBLtEzCrlsCrGsz3q+SUR+MMvZTo
eHYKFQ0s5l19lY3ifkYoZjtrWw8tjmJy9nWSSpuT6rZmZYbFKwl490f9De5Iqn7O9xCvU51q2SBT
HvO4aZ2CCp0BLg93lv0YgN/IGqX+OTrODetMe7uaONaE/ZWRQyq6g/gBsHtMJOZxafhwV/fIh3EO
ZlNYy5qaZqG1OJDaZ53JI4oaGMgsFFmAu+q1JCfEQ3o/jX99MGXyLBWdtkInEHoE46hxcV9e8lYC
obOkAGoBFIsxWKJK3Zm7EBiV823S75UYJAnoN/Lh64OLLr/50TzkD9rfNxnNXdwaopFmIqY7TZXq
oaodDOTbrX3F5saJrx5fj11Tm5kA5t9wp3nCrvtbIot3e2X9qxaZ0vX/W9xFVyQM4ma5LV3K5+ij
9HaRt1GqarLmV0pif55gEsKAedE8fbKGlq9CXt+jFk5YxYhCe7P9k6zmxgba7LRSNlVzymeqtF6M
T6gg4aGOZfxgDzZW26YY5DtLdaG2Oh8vyzDUoV7CrTaFms/Qk+5TOVLWZ7MR1Xv/pycUwOG7hkBb
izeNjC+qIgD1/sshuywNvUR1SSesFk4V6zdhOuaybQ5wpBJv4fCiCInswKYng6XRshJ//qpcdMb0
WigbC5AGF5STj7+klAwwTEJ5xMImQfUSJP0ULn/TYADWuHtfVPD14Ur2V7rejj2RIzD6i5ifQLsU
zmzaaWh2Wf6LkBeriqQ7PAs07FAVWwqUn+tGcolQw1mqmm1b4NFg7IYTsNl5Ethbs/zFLDwARGWQ
yKa9aetRXY5APar7ywcvr7LyEaA7P2l+NKlPgzfIfeYgltk8fOoNjIzooI6uX+gwQunXdmIdIDEU
jjZr2oGxONBpHRszdV5oAVcPtJOmMTxnoUX5KYWRu0pTFqWwCAM23Mm7W8G2W6cYzr4xcyxUCEci
38zssCBXk2roJ9GmOe6wPW8vbA3h8kBZYcjygwnwGEH4uk9GzLsMW6SyBMHLRM5nv6Zkvyy1+kG6
5lIq1BYpJzXBgVxpMVX1GG+N/ty1OY/PAmjr5cjxzBY9NNl+1z7na+IIcExQYlbOd8b0GTUOxztS
/5csMAmLV6x6McX1C39MjyLxADJIdq9k3gI1LT0SLRIb1vyrWc5En7he5QwFVD31na/VNFE16Mb6
Nmq2UH5USgP6kVqVDG1SRIcdNvO096fXvUwgQQJKeCCqqhR2pF5BW9uQRwtSb9ZhmrGnFx0z9AA3
drzDQVtjOlELOe4trRr2bjK55LKb4iXm8wqgmHI4g+j4fEWJVi6Ylx3FiKCcGTFD1And76UGrmyQ
1NoGCVJ/LQ6Mbr0+gUPZZRm4pT7Uvsesip+wncHH0amQwrk1/QETn7Dnbl6bFiXgl2ZQuBA1m2EP
+GSvTWt0nNc0uvtz0Bg9HwCEaHFQW9ccTJr1UJCLccKSZW5g/dw/BirHuvo7Er+IMDUy3DTFN9Qb
JfAAEPwXuQWBjn8mECz2MBmFSYWyJ6ryfknRLD94H5CKGMQ2fX6iZBPMuGgfYHnoYN3KQqXPn9PO
77NYyyF29BrAIPZG83juZxjUcNEQeRpnbREqDk0WeVnULCt9LnqvTAEur7Hf91KyjWvq6pdbYsYp
X1EFDMBomGB6Lyr4qbUxcNTyETQkdu/j5bgu815EdAJn27KBEnf+v7dNAHaTpbmzGjkTZsuYgfDJ
gRTXiy5P1c421doByYxaK6T+gEb2WOnOF7Yl2EBvdLSMLBcFNh6wbqKFRVpYgvGn+fB00RidI8ap
5/oSbqpJ9RYQazlSbWTG/66xwc3LcQ+fR2m1YiC5DoiBs6BdA21t82SU7/PdQLdtsBqSaIt/9Yk6
UFFJQH7w9cXEW5DkeRASIx1lIlth02Oq6IRaY0ljHxJ3zQsKpJYCnI+yIC5Uvm+XCXWxPfCauqJ0
fUOfUEgasNrA3ehgELiT5e1FuXMyfioji8egSFHvB4CZzV2FoTgpb/3cLP6zEIi/MA7v3oC8LVTc
aU9+PoygzA5BR57B+0nxABBEZj0OzCLk2VuYNCA1qaxsoKLgtcL7qGqCuMvyG48YPU52sgNVZBWF
17QhK6SPr4n6o/hnvKazNpJLx9XveEfqXV8Ict91hp2Ysvtz8qjmkdQ9NpZJh4fl2+jkhNxgXttL
28EgAmPvgSnJ4z8XkStAGAN50BtzmrmFodKakd5KKJwnicbkadeakmuBaGUgqq4gvaoD0uYfVMVS
Zr0M5WrY9+YK6vgq7VOYIfwrGebH41KE1+TYzRdeaeGdDqKJNivybtlyU5miV3faBzOtmn62T1Vx
jFHkAQMKFnIlFIsJ7S180OtShNc8Ro3H7wVFk/1FoKOFqYHQiuzLli7xVtOfL5wLZt1cmidiTxSD
IpKtAVHg/C6QbWU/0ks7wkIp0Fg1P/T718X51/Gd6oJMEbboUOdQcBWZWpSK9X7UjuOAlwk18OHO
blSrAXvsQ/+H/pjEcN4GEt7fOZdiw3KZc0aNop7eTJvyLHlLmROhO2Raki50VENGbetYFvKTWgaI
THzUxYKT9wOTxCX73sWNAkGqdgMsscGZgioc3gqOsbBlr0hjA9j4uJEQafJtDrfAk92Q+nl8ramh
NHL890liMBYZo5S+Yq3LyvqrSaVb8Ls8GyV5C2JQbnJnTfjWJvn1H0cmKQFstkVSj25etHSersMY
PjSj0sw7CEUrULYRrzayIUBrZlUqB8aThRISkZ1Oqmj9sKSuP5PlSnSYGVdrUnPkHpkJ4jbcUwN3
YEdo/QiMu6M0xux5CteqlEjg7440137UomgjmcT+oIp1kUjKXN3EXqKhD20bz5+QU/RixOCqrhQj
SWrot5rA1PkpBzJUGiupP5N5pglk+T+ucLTHBWPt2EYEBNVwvBuukoGkyNQP0MxXvSy6LmyZRDpl
WEYcDtjGJT4T4tkKf7bBlK6JKQBZ7o/e08P+YjY4hc4YUZs51qcPPqNVnC9LyrFIAVGZVyhoebEI
2wD27IU4zJ2jzrCtKSusX1c4sg3BbUudbK794WpWyekDl0/5yLtKYW1qMYyiTA3dW8ef4KgGIrrX
aEOFfcCB+aSgBn8uzF9TRBkJRtvx1ci4XWuJBH7yF7n3K4Wv4mgighgNwZ3ZxcNJ0CsLsjLpdGkL
eduGPRnpFLBTuBClxYRuYwtrw0KvBjhQ+qCqDc2A7YSR2j0xkrXSSb/X8L4XkzelseONmywgvauf
HoMd1GpJb0266q24eOBvSSfPvcClJBCwVZ3kFy0dAkkDpZpuIiQz7WZzae1X8TuHQNPxx8rjSpaC
biFMAcKvani6aKZmH1QKzhNIDCzgpa3rtGDQIaVoiykB120SWMqcji6o9ZfyBm97xjDJadfQ3htt
ORzWDWYDUxIpiVotx2tBpx/N8egRy7f7fwNjYCCrzl0ZLZ0H0ywYnd4P1lsRQs9uSX4j4HVPnkyw
52KxDALVyOQCYYrjHjysPT9MpmsdLcbMTpgKtioixJNZuKO8VAG6T48Yhzweo8eVOt6aJQU5cRTm
jBU6AJZe8/fPq1gKozqJsJrokLI3IOLqeKFE4y0s5XbY58LHCJ1SVsCC+vyzvqf1aw1dyp90eC0w
vbjfdI7kKojJMLZJaHY3bzfZA7aTTmPh8ghXbUoglLdKqXMPPhu+3vsYvUU2Dbz7Gbqgie/N2bcP
wbz3imVVLG6imucVdjJIwglKbz7F0pWbfuW9BBc2kIn2uGynSeYHg6k65AzJ0ejUtGdIi93bhKnv
1zp04fTtnVuRahrtaoWN4SV9UsVpx15p/0Ro9R+Ai2cXS08m3hAfZn21WdqZDotAU/F6+yvqZb0D
JzD3Ez17VY7cFLsxJLsui7xIaahAa2avIOIXOUo2mc11hOQTuaNL0AS2Ycc9D3yzegFcQggbiR9Q
DmjUmIEIo3TYh3jjW1qrWA210C8rBOuOZwmAErD9Wi0fdxcH1y0+FNbHueW6eNZiYGUSiW9lHUjL
iCKY/tKz1XS+8yd9RYNcrN+9jAsTNNEnliNg0sd9vXrAWgsHj/Xe86HXbNXqqUkBiV6Tm096+yDn
q+nxdeObJ73daM5JWW7QKm5bAUT7Wnd+/iZV+wJagrCJIT+6AileMu8r4Qiic1vwlbnXmG+s+kXx
ZxP7QKGLuD5lRiZ2T29S83gwLJa29og9pOdjHkBRfj7ivR2jXcs4h/u+XtTxsUOg3o0Lx0Yzj97t
M6emmADCogRL50BIsOa8FIfl6FAq61wbVXBbkMYG48bL4vVUnElSA7HM7coO6z25cvKl9A44AIbu
uaIMn7EXFqFw3UcrWyR+CXkslDSOyoA2OCHmaraxhss/yWFGr3PsJKkyeHnS8GwgeCQrsa0E6Xdo
ysGxZEtAfe4mJhmMoPcr2cACAPH9tX5DQrbNpVg3lvNMJ5ugwSD4Ee9OoZZeBLCstWY7NDJPksRs
11gBJywu2dJe3y74aaraTTRhxa+dwhnEHG6AqllH93wDg7+zqdKIywxcoVXy7GwvhsGdtcJe1XPz
3M0S83342kaPUdhTePOEz2dqJG828+rGT6QWclDg5td552aWroiiLJl3sVzZYTH02v6fqyoHZnt6
rwPUiboqhsL4MqTqWzJmFF3wo5qF5oHiVNNi1IzqCKAJ5WdUtCQu1a6OQw/ogUc1h2KDwY89fB+c
wNjJvG3sobpoElOnEzElDbu6W9Ysu/eg3++fB5/spxIM1Fe5/VezSExmRvepMkcGRMPSKKvSeUd4
Ck9G+rmIGFzp1YUy6lfEePY/YhgDEX6wcgK810DgGwo8r56aWfMw0HhKbNyn4JWacRKfhwyk2iqQ
s9DaMtJmwNLSbsODXOdMwqOBF1vfvqkiOfDdYF5FTtdgokbC87lAeBcB1XnS2q5MGR2k64x4q43N
fY4hy/7QXVovneH5mV/yrzOf2s5G4WIyeDBy6jcSdjLMMAY29+klFkDeTWNQG09qwhpBupRkMSrZ
3cKBUzL8U6n5NjaU5clOJhg+i9vDn5WfPxQd6aImcpU0JHsPYDGUYl2FQFeXrvWNB0rtAe5QCxhs
la8dJh3DQV/lTSK3wZyALoJiEf58987tn33StX8c1Mu9rXhnnQg867fpr75FSrGsPRz38LHHwGbC
fnkttQFK6Y/LX/T+iEwC0XnmHMCSIXdZ/n2V1ETW4EnYw+lpUB5QKj0p22+y3IwR4hwnuaP01ZnZ
bpbr0jU+v5V31ZJpP4Fw/ZIcvhgGBBWmQYqxoyK43s2xjx4LzshMR3hDIS8oBSqEj1EQxGoDXT/+
fb8pp3H1IXxF6jmVwcxRrB5iiMJhc/E4VdgzNdunb39GCGClR5utdHyAQ8F3WkrArb269UgsGQSy
9vRaSndBFOLMg2jxPcAx2kTzT+JuQJbWPeDTmbfYZ4exPi8Wom0ANaCLDOZLmoTgptVa+oOEDo5T
/wIlpQSONk/QTIiahcJPXCP9OBLF6ZrWMwDivTgCs+2h7A/bKliabwUcmVJGEwFRudNcsFmbb9Ul
Rd8M+c4HA/Rp2RKJJkiU6H+mlpcNW4N22BFzlIHn2gl8WiPlJ9CFf7pAlM6HgiaNIXyUA+0irhpd
eYRFDQ3cXP+ImSNpY8RHFMZ0PlCOO7jHY3UTsTZVxSJ8bUQThXuaPjlDs+z6ZrohAOMc6sHFmWn9
Pq0G/egdLTRdixSmvso73tNnWkhEccsHb2FmkChyPHmD0u+qjRaDPab4+yR3Vn5gGn1WfzVq72e2
bp4PI29ylPnxbV5maIf0Fl/1YDSVge6PqHJJNhySjUAHXzbYa2ru5YUUTtYcRIPEskcHMmR7WhJl
xpGcU1ohaM8vy4bxcY7cqoCWPKPCgKjHt+HxT9VMNYKJuIXe2/VRrge/6w2v4TQR9JiM6hZwoy6z
XGcayEQTsU26JOx6Nqwpj7Dc2xenifoh5H5w1k86cI7FM9cicwWJ7VxqmDvBpdix030SN5yYNErq
QP2Zc2xRjxDDRCGe9YgltlnIEgMbPKIYBXMHz6RmLVRJPmI4GUxIErL8Y3vCIqgPiPKJz/Rz5yUQ
7Rf9X8KTOpmNcQ9QVgvVFtFC9Pdu1LzpxzeMppK3BucJIRo6V5BvqvJW965uYI8/Jezq6nkfHsS9
4jC3QboKeVRsp3xy5VUFjq7SXGVFllLDrJ1JU8fh5JVZFMm3HLX2iMZhxFCAk4PyJOSdY0VjNzKv
mvilxwPowOZva5rHqqw/x+gXIeQNgAqkUgS8XqGMy252J3hZwDSeHAgpLkDXmTg9KlFXziTVQZvQ
YBpqCf5d3w+0sjXcwDeMg1/wiNglGU7r+YX2aOMBhGjfhdvg1GFw/qep/EvETxrKGIk32M6pQ8np
7lmFj3CIchgQZ7pz/lTCDqknkCF2JCy/MqvRJIhHDgCm1ASwd2owkl4+sun0SNtiV57pNhvoefMX
646H2/3IDNWnu0FcYQBuHKQSEKxeO0sCx5r0/8URK45TuEl1zZip2WsWYmql1KKRCCy90kgNzeZ4
3Ge1kiNR13l/kx4ZkX+DW9e4mZtNB9o/ZIpS+WyM7L7iCCEMzbtfIQH3bi65cGZIZ1tVCH5PoG1C
zNEslJwpgl4/MbAWRVSMJ9vnfJyCFfR0iBQhWNtEZjgL7Zp4hg6UACrhQE06AyoDGtHEkNTmAMDo
xTzrYTM6j5cc0zPDlzebzIrr3HjdzhI2EvOTr5SKSyqixDCsHEdoeJsyBkymTUdUVgMuZwOos611
4Kao5oKDYzYI8IbrXJWqBw9do1xvPI9ItR/AE5h7yBe7srKsC1nodpicBOsgtyBUEk3iCe4QTqc2
ubeiT80wlM/9dpDxXHQIqcqwdWxif4NaAFR7E5aHFh8lz9jgR3nZfcpEDLdjeW6Vf1hXxefi4U/p
y1xmupNOdwnewS+s+NfeIkIRjP+/odeJDQATHGuvXjD6Z7OUtaIg/KZkWyrZ/I/l0jIEld90l0EV
4OYqfip0yzrUTyZi1mPYyuw1JbivNNxao9m/ziraDkEpRyW0C5D3Ul4hgL7hWVtPdzdkUOD1n+OB
LGj6jAl6ZpzpgLA8QrEV+Xr+olJNorBFMNUENAYSkYzAdVRT89O1s/3upzY9eDdNh0elACQHLdZ/
baU0/P67ByU+J4C9l7tTgeQR+ldu/m2Tpoi/c0J0F5bgctjaIBfxpdZe4u0ALJXQUR5sXV1hOFKl
kg/iQQjU9rvxfXXqoXeV935xP9ZADdG1/iTfIAtUnoted7P8OuvZ1m5UfQfH3U5QLbxWSSxGqOuW
0Ipxc5raBae4erGJ0/z7da/Kj3f34a9ZzsFKbJFRntxvTc4p3imHtpVCCNWawLpqnYFrg7+hzmiw
zKQgry9Kap/dOZm3tQ+P19RM45v8grZ+HHmkzXGRL+PLohXTiZLUndwK2ngxwK66PtbWaTnzsOit
prcLcWbY4n2YvZoWiShp49Ua4KcvVqgj6CXmnMEyucADWEFARk9g9gJX+zvUhuu1LsdeelVFNplb
Zr7tgTHbVvVyjO/rnT1WzsJhm19k5nUKmt2VF69tgZVCSVA9OFVttcJtyJJ7rzn+6ofZLNmYFLeN
lZ1trcpRgLtkQ6rN9KN3gwVNs2IruCLSY8c4xkvNv7jbKmtdmmaKsJq0P6iOBsPMVmadolcrziVp
ciSJ/v5dwcn72IqPUUjD1FQX4Qnl8lp6iv870wXPySVIRZ7d8SW3gKvh7byxvL1F0XVOC7nEvar1
SFjyIJRPjoxnlu7ApyPWRBphuWcOaY8ImjfCt/6waNCoCwMFPiG1kDLJ7U1TQ3ShY/DB5Vhv5HQO
2/ZJ/EA71psGdVC4WWCO2SCBXG5+kfajhC3aStLOdLyJheCyBSuQe/MFse8p0gTedqmlVhyVk5Mo
qi8O0UxNFgih6ZDYB75DLRJ3vVUXPnrI51PsAZyUhfZ55JAv3jWX60VbsO6ZoFWcKVObJYAFEryj
lX2kZEifLpnKmsWpXxWAeYyo+pMUVuJPpIcvaHBsTWVu5Z3rv5f8QRDPD3XM3FYQhIuPcjzhT2iG
MgchhNzC5i4wX4tT8yyRAB+NS+JeXC3LWod76yinL1oFtD8oxbt+Ww1bbmghhBKcZenDRDReVGOD
GA8T6z50QyQLeqJ0FpzB/iuuXXUdrXDDYciV537oABObKWFlYpoHTHVfH4284zfb3g6Y8N4RRdSA
U38XwqhMD+U0gupjuvKQMF4/uPh2ulRZorbHRuoRjCC9WosygnwkqCbDGfvOMef3cJF8Nc59pYdi
DpqHJSmNxMFbDm4Z9u1aLV0ZESdMGUvzZ7xsBpLT2ckhTB6aEbs0KdCW7Mb3ZyVIqKg8WBHHlCrY
rm8InGJEHARH2HBAIXhagvwUUk8CAapufp0JS1wmr7EPswEhn5Bpi5NGIjTwopxkzqEzEH5+Rj5R
hkq+MvYc1B/yD3jny5F6MPtJdFcsXL7fB04Ih+C0j9IvK1mTGpSs3ugrGL8OrqPaJxCxfzVAsSeD
mGiFP/3nPwoEUhZfztArLU+Sm3i7C40GroSXkcCxMoJmngQk6tv9aZCz7Mg4Y4VbbRZX4xUI24UK
rg+u1ptf9hAodDOD28SOcXXE7X9K7ciTNQS0Gx8HCiGv7kuGdgGa1w2VNWv2Xw57zjytWZOO55YJ
USX+k6SjysrcUx3WCqFLp+/ku/OgW0Cz1XEtSJqqBXK38mY3Zq+0GAeVKNM7wfqYizS+Ixzg4nhI
GlMMgnG6dB6ogy2GGjjAT16gtq9Zmdgx5ClHHyawmMVVNfOwi3v822nJ+NeHrj9HC0yTuALzaFJE
TG+hrLmcBUvJGAcRzFKtxST7RDRHhz/BAAQBYIx6bp8VZXEwbiCFFY6g7PbyoXLhq6I5GsUqKcar
kZq4ekHK45rJyNQB4dX+5thjvWVVsRZjjk+yjn4se86jnwKGLts0ebb+u1DDij3gLaZNo9CwUMok
PL90y2G51HlunucT60pGmlGh3lsLCSDaQXo+5N3euGH/2ckkxQzf0cu/wgxhHc14fISSG3acCZuY
dECftIkBGDZ8dxU6fnue5NGXCrQHJyUAMh9HYUrTQzZqxKW72e6z0lN0YL7WyJc4si2WnNqgFNJt
aN4EV6gXV/bvl831RSFC4jjzLpxXlHlEaqfxttksj6z7VTuZdnxulsgCnHZlFkjmAK4pHyGEaOy3
sy+HzwbKCuWNr1KjlkYwYhGOO7dP3I7V5f+U3XHGGbXq6LMdrnCKWhudd0WNN+LbbF1MbSUlB9gm
/HliYpqrtwEFXCgOenGMwhr5TaTQSsO8D5czR54M3Ai5qTTSdkS+V8q/3V8a7uCkrnttg91OGjEw
sSIBBwbuJG6Q0WS7BvqXZUZDHdDn0q2FwHziNEaOycuQRYxqAGWLAupYu9KHXT+LE9owehFHFRH3
qpUSgsL6+BQNoB2bCs9P041S2pV0zKuoTxI1JIaaQGfWCFNkLpY5bOrnl4pIs/TRr7jsJT4JM0O4
PHsPOtJWC/VSW9L7MJYbTJO4pyn/hCsgkLVzd0O4nNim9evlWab/fk6DjSFc6TuAIj8eWLkWpye9
m7dRY1k9WQDRdf7dw7YM7Ig2C0oLTZPLs7TihkXO9LQaAbMVwnXjVpwqqQEOqWknGiAyEopQqqBm
AAHJ6AONaUv085CXdIbXQ6ENHfp8gZToa0E5IPz3/vuDWwDxaDzodFlY5UE/vTEcCafzPgq6UvKU
QiOb2C9o3v4l6I2o0QomVd9wlhH9OYB8gaaxavCCbSKWY5V3R/OGomkwKu5SsbAygLPR3nZWouX9
Yp+58xoOOGRDc8gjENrBHX0x4eEOUJ4AJl9SQZmO2xlg0ea6P2MSPGS5p5PQqFuFibKC2r7nTEsm
/ij7M7YPhBObjqDfFSYz8YjloOHAXRWFP78Pffs7idas5pWhgHG/85fT3b8X+6HeR0CnVYoYT38E
DBZ+R0ibWWPHvVYdzYyKcajpnd5bhfXGw2Xtg/cPf/m4lgPhj09UlPH5YoV5vKw/WLy5rcqDG00F
YBvsmuBh2ulf50G2feoeZCy5fxDwqcIUTuvw536q2tepWeK0D5pcowAi6DqWcWC0BXvkG7Xqj2zQ
BXKWg2AsJa9sQyqRxuCTeSgQ5Fl9//H41sm739CfjduM1pwhtSQlG+tiCbnSlDByiK2urWNUIojB
iOCOzrgK5i+Tn9N9W/igwJJWhV0Fg7sEkbDXwoiRlS2Z6TI8XWWJ05ignjjBZHvj0cHAAHDZNJcz
W9lcEVIWFFP+JOi+T7BU4Q3+yk8rQef0NPuzw8n/TS3QLYH7Z7KoxEHcmIbKcAoUKUdUAeaWmuqL
VG757UjVX5zTRLbsNy6Q8PfsDD5QP69eEyp0a8dtLDXb+gw/bg96Yt0ovcGvON3tBZxbQ2M+jeWQ
hBmDHP+3dUIFFKWBP5OVeAYxNVo/qOQrxRwrtIy0MdlvDsMf7jy0IgDwyYyFt94kc3OBU7UgEJaj
FRl7hsZvicdxWjjI1VHj4IlP33Tm1M2AifeIQjlfEMKdoWJjYWFdNRLMXhvhm6d4FHfY8b0/N9hw
vo1bvE/NNIWlEo2TZq732rKoiFVcrsyP9xEst6yAzqLWHEjw2kjt2vjoM4p9TOP9ii0JBYBe63AA
9DR+cHPqqfUMB/4BAu+NP7iq4yijd3TV/4Y387yWScXRpjwxXwsXvREjpAVMuW0gbcHVswvluurZ
hDiNGENAaBoscldoEJDXVMTAupgqbb8/bX6+7xUIzZN/FKTJPY7uGLHX5mBA67VQDrbpLt48Aif8
yiK8o9Gbp3wcewdXHxuuU/pE+tkVKZtKW8ihAOkKCntjpHQuKLw0AMJkpZ8wcN3GKhaWoD4gry+z
37snWmqVj2Lox+fzbyrzh8JbGAVhX00in+G4KDeC1wwDqY+h93Dd7QLKDKJrcgbPqWXzEMtW8PWB
hImlmGrbbHykzYAh2Sga0olmfr4CjjOmlw4mAErTlujfRYunV2NxF7FtZEteUJkUTCvzvAkEG9ra
9b46h1zSWtoLFDyic9ZT01YKe4ebggYf22pteZFxkaS/kYCWvRweHmUYLAALwHFy8pRyseP6d0+D
WBoPMDM4BPz877OnwP3rYKcF5N7O3OazZR0bAE7kqNxs0AOZncx4GRf/lw9+5DvW5RPUp6FpH1vp
kgjU5wnPkfS0/MQkMIhQh1z1/leiZfkP0tMK3WNOmIPHTPcjhJhsNXMFA8qGSyo+Pn/EbH1kVZDB
/tBFX5jB7ByS57++lsGAtw5N5YJUlUOlRFOtULK/3q9LzlaW68lQ6SnfRNMHiIwQktjsGjoMaT9e
Xdg9eRUWDK/1HIBXlAy880p6RbBCc4fG1FqWoYzu6Gxoh7xpfWwtj1+gAFZ1yxLKTgEs+0MiKIkS
yugf5JGn9sIxgKZ2U1KlM4Z8vnhRpPW5NUZd8vkuIFKS1jbQUkO5x3CuJbbPKHVxiBJi8tfCqGC4
pExQ4kpk6DuRg/kAsyfXqxtW2Yp+dir/IQLhwk7QSDYCVbPwwCF6F94TvUeNP8jP3pNriKd2W4ms
5l6gRzRrQ8gtyFScO+3LF//Z4JYAwz6Te7O82N1yIrs8JK23vTkL7yXuPYiBmHnyPndloBILfdqZ
czpTCMZO+bUP5qw7QayfEG705FdFZb8ZQbpMzWfDLM+Xp0VN7aIJWQqUpnRTtGabbkDa0hEZwuUv
9uQQ13XVvLeEQ2l7V/XroJu19ZqCCftiGMHqUe1mW1y7eQElohJ/KAmA/MKSXEq+jnQUM4TUcNcQ
rT1ACJqbalXhq5G1fkpdGc3UWswtDDYFW08lshkjOkvRk7rk+eXosmfh9raI7JBQ4O+FmImNkrFW
Vi9rZnkoKbLddWfrw9Z8QeptaLCBijuUHEzMluMGlDnrSEowyyCKdOrg3XC8bWYkDP2bjXaUUTPY
i8HvRKSQ801t0fVPYIaz0/fVAg1M1lp9slgQlC9mU+gWcmA4xrbugudxj8r/4vqhCEg72lE2KeMU
kloMCG9sl5chMkFW8luodKketgzFmtkBfelcwklHjC3a0HkjW//JY3HlBgP3c27SCXrCTxAwUDs3
pQK51dxo8otY9a2nwYdkuYWYSUA+Q4w99OVa6fi9E08SPvF35lSQWF3yQlPV0ovUUc4+pr2fs2v/
YzNwHqRrK39R+oN//1XFdLPgfMgCdiuCaAHr5Vn1Qz7aYIODa3gUoF0ykFUFVLrBY9MgwuQwurhm
m1S0E7rJpGm+BE6TYNVfHEef0yQwrzfn3HkgEYtAFSP7R9tiXAPgwZ+bDx7XlhvTkK6bmu24Wbwt
fZmu8tP0DFOD01jwlJiuIDmqe6qC6M0zsgtFxH2emltptLOM1B1M8CWksUmDBwAJE8K8D+t7Jn4E
Hr3kj95Cza0OfRL0ES0//MeBrhr1pae3urkU4ZF/Ne/xPnWEp3bH9UBqLEkcX61Q47psMWO6NDJW
d6LUiD3BL0d+AFA/FDIOgRt5eUTdvb+OyJKhjWeyCv66BSs+sSudpYeH/aHtOOMDU/oyD0sp+fSm
qgIurXGocymb+Wxto7Qode9OfLprjJAilveElj6B2sqbxttWSD06cfjlKOxyuw+jf1ZQK+oTcPpW
R3+bb9FhW/9XRHf2H5zCNHVWKtbF1O8Hprsvo+5JoRqlggLzN8M9YklEMwkmeMNuedtmBbm8lEg/
VwfNbndpj0aF2Vaag/rhTf3z4tYBhyAP4xtrlkkZ2m0mKTahCpz8eKe3BpMW7Yyuf+hnJFParDMN
/9UgVLUG9tlMljpm9mIcj38kauR5K37mTuOGwqLU4DgIqs2IZRQn2vH/Vy5ry4QdFhynoFwt33M4
AXSgil948NJrclZF7K3BMojhpMkUWXD4Bqs/AvLuLraAyefovvKCmv/+6aoTIGgyjHAxR7PWMhxc
eermIfugEEsKLvJjhVUyUrUQIr1NnTxyfDoqUxhwJ+oECPnDu4x1OfdbNhS3/DUJhFZ9OTYw6cwA
3/I+yo1jTWkgCv7CnOvzm/Hxt+2ceYr0bcSxxoofoNae6slO6IY748GmPe7O/4dQ1kdp8LO/AAMV
Kjj7ELQVMez0LM0zQ2iNngnBOTLZ6kC+AjEHLXjCZ4m7zHGFzk4cbVPAmL4gxDYPIT1ms/W89Ewd
bXDkdj9R9cg6uRL5KNR/1KHKcjyujL4CuB6LIxs6NFy4gDbKdFWP/x3IhKEBHFudWgfv/0M+yHF+
bsil0CX2SPuAieqis2NLgXMMON+4opFBcmRjhs/aPpyCGq/Hjoz6O79kD0rYd1vqGbQ8XTbLn1SS
EBnjaIi/pO6N0YOwstigSNZiH3wMwhxTksOc0Rst42kig3JdXKpgH64y/ymHkhJxDOHLsuR4625n
fSLZ16y/vCbi5ASUcpOYVrDbgLD3FpxVja8RF09V7Bfr5VenOFDrXKaaa4/QKvCINXlm6R5Hxcs5
3rLRBX8hjNFxWX2LYrE4jL6DCrULdcnCeh9O1/mtzbb7WG8Mcs3o9AqUVFN3xJvPg2hlqeEBpmtN
cPmSFoMF49pswav8r/e/hIK/+aoy0XEcwiKwVE537MnsBzV4Tjv/tuvOD2M0W7mvnvTpIvIRhfEO
G4c5PfF2Uzi1qOkuV+wM/Z8kqICsqVilRmmsiHDWNn6+9aWmEGs/i1KGPm3xA6hvllTv2fuIYoer
SA16/DPjgya8FqAmUrC8JH1BaPXQaWiLdbYwV5mCE09EifZgRxJwbIalicyzfO4YSVlu2YAaRBWC
dYPe/+4NkQFKn3eomMj7exnBbkQqn7vpv8ldELIoBGBlyAEt9HUoFa35lbN79vtIQ3HpYJt+jZjI
QdG31GAnmbmyr5UJtltNplcmn6Ig+UpFS3aXb3u4VB50xb+nHyD+c0wGSnbBhWjL7rKKeGIMfQWS
8DaTa7SFZinT2/raz6K9vxPsy9CIDoM+8rDSCWD6NmY16nqa+A9SWJe2OkgPlSySE45Pq4igGPbn
0bB0Noe2VDirD/tLmWkvVLOnWIzsJtz42O9xIkmLScWofczv9FHXH+R6q/9lNQWuZw/q6p3AyHpd
EXZz28Oy0e/D0CeUjFMaiU1Gj+Ex3zhalwKAs6u/j37Bavoe3SARmGSbP0iqG0vqaaEyY0T0aTtt
fbJw7CEdn3yndKsyjme/9bBXD8xyKnssSLxcynCRTbjv2KIwVnlj5Cen0P74cpG7ASs6IIaG66fW
gMvenvEaCqPABNzsaDq1GZln/+YY8Lxm2I5DUzcEAUGhHoMZGgVieF1YW3DsF6BwNdWVQ4mGFoSp
EbMXVVwN1qQQS+XwvjkwN5cWeWswHtJYsY6mHHG65OSruRGZ9OuabU/64v0tnA7v6l8B325yQrvJ
GTJPyO9NLuTSgwGKlxNpEdkuX/lq8u2UQ2DbrTohuGcOTTQh1tctLs9he2UBNZpcy3LgFi94tpBT
HSjj3PTGrEIPckO/X/msQjWEkkLdx+s25FhjRdn+Q2uXFXAI6vV65WUduYfs2DO6yPV4ufaHFZEB
jwjH0GvM/wm0B9zOFQR+bLhwrg42/oxzw9QVjEsRZhM4220d3nWsnm+J7wlgK5obEurZsc9zH6cf
mDylp7uY35Y2YAGdlGXI0d4VLjLI7KulsBz6wONkOXs7IhoM+yeC7o9/vQoeJve++otRCgaLQvOF
rgeRGLaoIg0EA0/3KUqLE5ucV4PJlm3jwu+D/7zHY0He6uyyQ78vihRwjgaswWytnM08Gbj3NwZV
XFft6nmPFQ7M19fpW9rGrYH43UijNbDF/3zCW3G1hZ/GMZ6hRrRc3K69sapWXBc0Z/B2mvh0k3Xf
+dNZY8vuUTJ+ta9Fg7BS94h+Ghj+V9Y1Img6xuGqcKpbR2HIJtR/1DaPc7ozQfH58RYTLupWlFAh
utblGL9WVy6Am8apTS1Lm9+q26slGY9KFGfPZGm2I8KVo0q1asi1VQMCQGYhcUDvsWzag2b/j7Pc
pcdBEgC5inYAp9L/27OdfdZQ454vFeUCqJ4vT851F9EWtety75127pzxulVDLoomoJ48JILLR9iU
QLjjX2SX//O0FAC+uP3grQOtOyErD/NaZQRIgesFD4BjjixkN8zrdjMv7na7AHWOTl8O4rYYVDTE
Xql0AULLUhZOqqytkyoLpVUcLPBF61+TtdusLHJxJuMDQ+DOaEHuxVaKK+urxPYrhrYV781voqd9
08rr6hFv2Bmlw3nd2AbUjdus7T24fJZjSiFbYjYqYKLnM/knq4lKRTLE5TRJsCaesJHvzAtUwpLX
OSH655VxPu4YsIe8CMQFKqxw0ud2Atl9XSwAwLRLjRWO2UJE3dGB2Ky3To3bnjJMFSilXceeX7gk
Zd4hpQ3Pf1HlUuKo7ehfjQpDtiH58IGkAztVhlHbNJ//B04CWdulV8ki8C85r3D+hJjKDSK4mwgO
0xzhf0MtBJ1rSX90ILofYGDOGFDcWlokBvK9gsBYB7hUoRnPO0FcFnTE4ZEERXgy9QMKPWveaWI0
ydk7f+mqzHbYSJZtv6GbCN+Vve+SJgOoQthAltDlpK+uiMKDkOAC5VyxTeTANGPNmyhqoCl6V15v
wjMYTNeE3ROLnI+MKvoZYPqns2Qo5n7uQ2zPwwZWukKbqU+9381Lgm8etu95VlnWZatti3NGY3nc
T21VnXrq3v4QEvC/5QXVniCzUgt7gVujZiOxt0ms3+aWwYSoxtGXEUPkjwqMmdnbPfSGWRJ5ala9
eyPVB9oyjxnq9hvzHFStWjpVEdMO3CRDcGXICkNEKZY+irPIfba8ii7+VkG/Nw/nbz9YSNkePGE3
lpyzDwccSiZlATp0IU4ltxtTZ6874Y2aeXsi0cZ0G6N2tasafHM5f0OCUHd2zxrpDJtQz+05lFPZ
MvUXmIg5InLTQ5gB3pyzz5yclmoiYGIIJp1C8BphDpbqRWqwHXrjYgS0QLvOOf91ZI90dTo50yaK
9Z856MJT1/6G/S9D+gXC9YD5lY2wDON4Y6PYSBLMAVm7MRGdBwbD+3q8FtmIOtgDpczlFYoq1XJW
seVClQ09jxqnb5I2KwHzZ89WKe6yc7PMVrQSxoJk1vNrINvR3A/eu3x5NNOCwd1MUDxgXcO0siVd
LLD9vBdZDCJFnthNUukZr4PCE+9w8SS9IGY1D/IW78mpPTC+hpUsPHmGUTd9TdkXvAd1YCMxHXQg
FGMv0jy/kwgo3bHViq9XIkJXWg0huLQwiw+tXwNOr/1THIz0x1TmrRdzOn8LanClg4Pjn4KjPuIK
TvBmYIlIzGqxsbTabpvYjKIBwRx7sSRnoBGTAGIIROrNMs+YSAhy2HmsvMOg6wc0yBOuPccRPbYs
oaC5N2UUcmFmYTzuOjiqu/KCB/aIx5kq0B1dZ3RaxB42essmFlhqryXZCz8OqaLaaATQT4SeEu8i
FudxFhI6J3iYoBioxNZI+yxhvzG1r38fx/0QaZ5Syv1n851DzXvRGxgyr+GeZS1FFowzTmkIJQhc
6OstRT0j49E2AFuApkIeb99sWnrHOKY7sgqMKDClgr/PQrRxNO+ACpTBzraz+U1V+NwVXqyJoneE
3PJubk9b4tH+8hXtWlWm4wpSVTecm5FRitpYPTCqOdk3K4+ZfsfFy5y8zEEaVUh4iwWYcb/TnfTq
9vuEIWuY7ExaRZOPZMG+6IY+ptK5qua/KlGccYp56xS/Wo2reRzoRJOeeuqqlTrDbGUq5HIHY0zo
SxtHwzSSbxPANAubOG/e+xinspb75kmrVUqLwO3qXURQZeN1xdeA/gLgjz7VyKE+/tu58kqo5af8
p5vfNbC+c6MagTGrS+PQzbxO5i6CrunXgIlTBXddZX+acKc+VsMdSN0VopZVA9y3CqJaoZN55A3D
Npjj5VbLQSQlbHeu7xO94t+iTvlAlx5xHTJ75i0Sae1n3TuqEM+pgMLJ9izGqDHmAn0ASLJ9w1AK
wJMi9tN1WI4rbhMugLWvXwgoJIkMttN6cT/GQjJ7BRLsxCf6j6fsgs+4qXiXqx2CvJ3IZ30SOEzO
1xxV8mohJjvAozyhhRkByDFvyo4GjqwDWm5MedP6HjcXomD6RviWUToX1YszQ180lPVHz4Rn6Bex
k1/SiNjnD1/h0JxTPHuhnDy1EaQbLNhKTD+bFh6rcJ5gF9XDkoPPqk1Xw65zKiC6V5zk9De3iQlS
BGxughIV5ytfQubrrlRE8IxjYYj0TBBBU1Q4i9HSO+9VOHCSdRl5YY73yvqfwSaZTfhIFqAofSIV
s8hRl43Z2wLA0Il8md81SX7F7haf0bXAQgzMWaD6mKOudXOu70reLpemop6scn43rqnnTu6VV5Mt
lVE3DI1RZlYZ3oAyBNKWDyWMeCG6Z5JsO8+19b2/xMbIEWjBYX519Mtc49CHxS5diUqOB7CZQjKy
kbjgk6Q1K4MENpX3CC4XPSLZHuu3JONLElNuznJSu5TlZ/+gOp01k8q9vpGrC1qjJ76Ylzb+Drhc
jrd9HKjbyLJbwjj2GulmgFpQrrL5VXG8wNNQPPAZS7HeElZv92bOHrwsBU0cq5+kuuAqqgdRE5s4
WrW3827OOrMKX8jJsW9C+Pz97VfGFi5/Xa3LPcqAaMdn8mFjOe6PRwnOvWrGKqkQNKUETD8nzJcm
UsDB9IRBg8c7uJydUjy1s38uvgx9qn7q2q7HrXXP2YN6IbU9eJMuJlxq1o2EEnN8uNEhI2i+HPu3
KGmiEaR16/jrGl3SOrrE2AzU/e9I0LZwCokunvqbWMXpnyCgTAALnugBFufbcooPi/VagQnPur8p
o48Uf1y/lcIVqtTlDmoFDr5AFv0eGvnT3b1QywtcFZlGdn/beyG5dKwtn/cy2ZeNsuqO0vxWqPyG
fN27ybp7jp43Pwf4WT4YeNTkcyeYvZfxeD2IuwW21nKYqDZDNA55iAHUZp0qFisqqZAfKntYbRyg
4jrhecQDMIU67eNZ4vifgEHfGyKaDXF5r2zy9JBP/S9GhYOZdbqPeXrizGFh0tulYvtczxZZ6XkH
Z7fgH+tuyC7ovtdycQLSzWPSHlMZVrJcH6ET8rgahJuIC0hBsagAiRCv74rSnJKwcGXI2IJAYtVm
xxfAWQuGXCf/mg3/msklskyTizXYg1qnGfMBFhZlqnMzJ3iAp8qYBJkL4H9WVzv1BuNtUablnWKQ
3YLczAxfx0GnKdq0GxjA7E6bneMO3QTg0K4UPXfjvgxO9juq+ycm+1tstyp2AkFJ1obYROVi37s3
P2BVSZUeCLchh32kPnPvAbar63HW/y6/gpeF1k+yulRgigK0w9WbPIkNV3OghoIWRzee/DYOcWWQ
a/O3HTkNBlck04D74EE6o2me/Gms5tqpXCJxF+ejUTVpj1lppV62OTXOia4IgvW1UNO+2ag1fF1M
PCj3vJVIjMcVzMqdJGXhPYnIZYCozgQyxNdWhMErl7+pHrqxoZx80xqozPqI6I4UOV9ocq9FE7JM
ShyJ3DIUjc9Sxc25NTeqrF2f+y8Vbdg67Q/dcR1/x9SvrN/aZ5MRuNo09buIK4NyyU8OempkPDNa
Lh4QinG5xBx/rREDknhcI9bof4rwm77COD3Vv2003to6898n/QWyJnBYYP/vaqdvKOWYP8ATUqiv
0Cv8p4qHkvSbnljxeIjC9DY3m738brXmkRms0yiNxoQYHDACN20z8mGCm/ZKLJLiz9Dv0categAR
cwRkt98v8jDBazX86rcRXEEwQuiSAusA4lWryvMDnq65mID4B1WfXLom4BWthrAc9/9h7O1uzUn+
agJsS6diq+KrYf1kd/Nt3OfFguXWbLgXuVkQb0MJ1MSl2eMkSY0n4PzwG6Ev7TaMN+mDF2Ohkr1i
t4gr03hOacVy6x3LhnFExRiK2MpyzIsECLlwiVLub64OAkTikZb6z6MBGavGeWbpPi78vMauLnn5
3cKqObW2Uv41cYPKz9WcqEBjZY0AAy591DKFUNNJeaaW0+FPjj4IpkWYPW5VGAH4r3lCs2P/dt2u
vpllVuOz58fCQ7eUcxX4DQ0EQT6QpomhqrdieLxIXScLPj2tGmDpiuwk3+zrS4zCCIsQmnw4vkrW
DQLIdWm4KY3mnuYaIqshgC3/qtSjFNf9TmXlbSc8QaEsOwfkW6SV0aBuqNRspnfKiYhngrNirgAi
rPlyPCZpp2DObCFLenv9Nm/Uos0bqM4xT2+VEr7mqLJYQme/2MwlmrP43wVgMM7H9hmDqruURk88
++JQO1Ce8gLisZE+BmFZXLdnrUaxl/tAt/zwz1nQx/zEEXPyTsqfiveM+JbBpBc0wHW+3YcKmkFW
g1hkO8vXMTddOesDYeF29F8JqajQn5MW3itBMpmolWzc8XzXTS/V1pXuYd7kdiCJ/BKBt9iZvLWr
vzcvVSXnShlJxjNc4k3CU6jbCpU/r0QlJNwmMUqevP+AHDDe0Rv5cLiwh1qWmz0JxxNFLZlkh9g9
Ucl/nUNYTMldMDHZ1Yeim0Cj9SBSricC41k8JqqfElVK30xPoDWrQ0lvO6Mas7Q8yVPt5dn91B0y
GOONvf/nOAMoT4D52VgGynYNN5ErG1MjpfA0c/xXr/t+5fDbvkIIwKQyYjdkBmln0YFzN/Uhmb4F
kuA519F5unn8nbuw1iZz0B8MtuO+SsEzWnttnzOaiCg1bbK+msOSLY1hi7NSFlChxU0YD/JC5trr
lpMtWRAhxzDYbO1NK82vALGF+B9qV3zpZ5MndXMfJcFSyBqp7GlKF8JsHoX21ALBWW0xWot5YCbx
ZjX6y423RPX6DESrJTx4e+H5MoPD7YwW5I4ZmE4nnb7i0HliFaE55uZsKd4EUy7FIzdbdgQOHMJa
PUsawxOugd2JgsU+fuwQEjBd6/qPbpj06siOOHqoMk+AIVyK0InE+ndF2qGEEOVvdVXWxSjUWvm5
EL61XRAKTAo5DOPGxs9XU5EtP6Y+7NzqYzm4Htg8Xb07dx8upAvr9DN5Lu0RIp33SFMWsefwcJB8
fN7cD0keXma/DOGH10Sbc3si2VVp7fPKlZmQ43aaxoEMIZK8RPcp7GWWKR5iPMM0Y78Ot9T9DcLh
OvoCQqka0YyyInXc7v1+pZH9H2w7XjTrtM9JrBtx7ETsgk3SoZJf62j0e73L6WTfCAEr0X1M7izP
yWcqoGi8xmia+pQ4Jvn0C4Qd3NAJN6tV5FORcKoncz/tV6Vk1ffE7sY8QV+emnis99COEJL8ihd9
Kb21JaITlVkqjiZfyU4Qp+KYHeDLpW8UhdbceK/D8b6LZuV5pZZGX+lVtc96QPuudJsmbyiLzBwM
EKiEmtT6eeEq4qnq5bNqqWvUHy9+D7AMkp3ho06JYd/WbqRg5zav/+DotMQ6OzFnVhQkrkbDLA/b
qNwylBS8W3mgrs5OWLZshl/dH3tAtv+31k22pBgNvIyDCSw6l5Hayrwt2RVZyhWZvnw7nlHAI1bh
VmcSx6BYyhYH4Mv0eq7zHhJGOrB3usouEwFjFOorXmXXa3JoTiOu87HrnRpQC+lcb9LZ9NoCq7i1
RCQprPXDxgaCXi/RvmoP3OK9lSbz2Z2Pep86rHpEUfCjieekQcJo9jAT2YrbOK650dWQ+y/oxcuB
EOll4vsoqPrYvFIoBnL0McIusRLpyeQP4HARfUcXqCKCQ8viOmvNXFwTO75AQe9sV/u9ONcRH+gF
6NtSxIlD+hqxqzYQmjhn3mxDp1dFs2tT5kXECjEwdGbtIzHS6SfwbNgrpGKqtZtd5NfGWWrrLf4C
rvpaVwDyzNKysd2HYXraNNaPBNTcc8s5O25c5J1i0FJTl2A794ChEz6Ixxp2AbbrzwEYhzw48Mw+
PGxo2PvFPY4jRTjYNTs2ni+6yGzvoXLslACBAih1nsZJJ3nKrbLmOKzX7cvSLvDIpa0+UC4WtF0g
zPsJ1E28DlOwHRwMfROWFYNovqSH2vnBvRPBksM4tSCg0RrM9rgcjkB/S4Y/QjhCRgPH7TWm3Ud+
zl34BNmdA7pRAtOIqPnj2Do/f9FKf4dv4jkm4serhXNG/InbBGCTdXqp5N9c4NorD2VoDpTBxGtz
VmP6LvbIDDTrPDj/Vk1B2d//OTERvHZsNGvA2xjuDvxquR6uZNztho2dLoirQEntnulSbS+BJ2iW
upCcCLORQxVMx3WNSnEHAU6wmpbbBO1+DnLQtL/Kg3FfarqBeMSPJETewuz7bKZnUGzyuwTBmtC0
o8xZWpknzseBCO8TVAqALdpr/5P1i2Shykyrj0zhVy9sMosGpe0cu7oimV9W+39d+LiIPLuhj4ju
6JvlpqRU4ysmdaoowwzR09Vahj/qSAEW+1QYal7qs29HiPm2i2QnJmgOLalleq0W38OocHwLfaOA
GoJGlazbHOEmDhca/zhXkc8bf0E8bUZKwqttrxq5W4QXmJ4KA7JAtS5qHhC5BxCHLrweBmku3vol
3VMaKNtmAT91Aq5nj1vdo2JG7DIk9xIrlZmonYRY6xFx1Ttmdwqbiv3xgae0R74JiZ+J5m8k00cb
lVIRpfA1SZ0vyEkScO50k/LZDAj/FlRjDsSTk8DfICI5l/wo+k7pL51hB5E8i4vVdEQ9hj6xlZlZ
+oHVZI4A7RVWbnxSvzDZvWq6hadRD/4+Govbm2bC01/GzQZ7rKchvMjH1NU+F/qrIEXr+N52tP2s
otxsK8fxDZ9FNit8lP/wX4JjBRGwtQdU8feJFYwa+pGa7cEVmvJ6S5yYnb3u2H71Spu3M0ktyl5r
6AqH9jm/y+YkBU3+/wYmHcQTCbHR/brGX4+GMY7CNBj+leveieOV/u3gjmkVSGimqk4AhiQukgP/
dAgZjJ0B4+9CFXfcVKvW/ofxyAt+xth8BUu87dF3ESvyF/eXgnGmOAZVs5JMhNzwKzp7GhuL9r8u
TtOquZ8jjp3AcuDwjSaHuymWHbyc+pmc441kbuW4MqEelsjywO4jde3vjlDyC+S0lSLGxL+HFR3x
6o3kTIuCN69huie468tV0rrhKJZl035poPtsUt6pB9KXaZ5LLRYkwOLIgwopEEdvVWWSKDkMSJ6G
LCin6Edot4v2FHa2RkSEAK0toqe3KxJIoSL+5k01dUYAmK4bESjZRSYNosi40g4sGWKK4pioJF3o
hiIrBQtf1DM4+qtjshZ6XpPfrJKTuFDGq1E3mb3ws0dxGo7LUH6+ORgP+4OM3JLpw2QFIWVrlZAM
6hTAsYny+75k4nlu+SaAFb2O3Zt/UuJo7/aH7YTsyUMQS/wGI7lcDZ3lKdywZx+J7i+2HZzUJF2A
POLBT8oOWwrPvmDdu5Kn8QvUsCWOWXhP4U2l7GiSweHfZ2BUBOxy0OE8QWeU2C0xdNWW4ep7swd+
UAegt4VMJPcDG5so7Fe3h1jFXkowDSBypUTqjDAj+7wbuEtGREMMuZyv6rXcGTS686Dy9pcWO17R
2IgOvSAQn5VRTxtGTF6Acx4l+FkYQ/LqrnwTPpywPcEs00GH28S5GBwJ9yeZze1Mhemv6xwoDsbF
y+8x3lJyW/mZueOd70ExjLLQk/468q7zy5d1JHc3Y7HzMIIGln2zeQ530/20M2bNLjQ21IjzAds4
gXmkaQeRzuW6O6EmQkxBCwnzb7IEdNwOyX9fEY4vs/vyYEBnZgJETABdtqasF29y9BOkFxeXsnZH
Y5aYMuiIp9rsmxOSCAxByyO+C6sUGtaIkbVWAEaz0Uor8Zw6AF7wv7Kfmu7F6WL62yNdAjc+/Jtj
HbEc7o3Al3SymqRs4pQ5SFdcI6kptN3WL1MCaYNTYmwwTZF61WJ1nazYCTZIGah1mfI7zByMHjed
8fdbsCRsOaHrRGKblqjegOsgaaSxUHasYhOHXOgM8oTwCHB8e47WI/HFH/tdNv21zLp2P7CJCBRR
SeK4v9IJp43NiVqDxexH/VDjzRshrmjLMFKTLBOlgYGNFpV89qUIns4vW7HwdkNOqDZmshi2xiyU
diHGC1ocF/xVixCfqX56trOkcN1Yw6WlgCm8A7ATP8wNESgRgnzeEgWidOx2gxrOfd9H13GEYu9G
b8H0QUwzORXkORbmmeqIz16/bdUSBA2CRVi7GuSh2YGfCGuhk+JuD3CIqOkwLHpHEH51qHLW4Wbf
RJUCWRQyvbTnkcaOHJ+n04msG8D5HsQeUGx2/3pGF+jM4LSpj5gg09WXJvUB3h9pog8yipbCOzFq
LWEROitcGWfI1w95K7FJATaiHX+BVQmiHxvfyhU8PHJckBPtME7qnKV1RVylMpDVxMjUhOVKB4uv
BthxlkHwpn50l6sWPD98+PHPx4/qXaqLp7J90Zqp4mNTUjTgEIvffgfUV/WAbiNRXAuBBqYbJrTZ
/JNJ3M8MviizT7O1rHfkQXWXV02x7S/e0P3F9GBbMMq3CJbZo28VpWbtKeJNveELQoiIc7vC+GRd
bMbg86WbEDnHVy4ZFyjbcCm+fmg5W9d5WlekZ9GdtbjHNIOo3rkC5RdllyCXIGFGubR8wKUavQJU
2Hol8G5Mu5jYen/BBMwUZSdGjNnLCYZoNq20pW4byNMVi9LkYJ2tGjrMYdg0ieB6M90tePxjVdwc
Ib+s4E2Honq9I71sSLAMh1P3Nqq5FcdF2LhJ/bKKdBoOH3VuGVjBw4lGCK9thBwqQ2ZI32OlZGo+
wYBF+G5zzioaEWZLaQDGnLg9mt/e3YQI49pCeyd4g23IxYJv6PGbTw2R1YtWnorzOISn08m6e0Be
FDMmgAmyOJUy8UHCDrogqfEHKGgxJ3t9uZi+Gt25DuGryQ+DWhA8p03RcWbPS4o2Re+qmJDP1dtm
i3Uq1/rJvltLsTtOwMyssQqfjIm0ssx3KEsUyy16f2w9JwCQEnA9kQkQJziHzt7lzHMo1UisAJk1
pup9x5wAJNdFS1yEeRfvAEYmPyg3Q5Tdnyk23eIzVFruD6aCtCmlxQty9q6/xmwT4JUq7K1UrrM7
VPWD/NiMJGQx+0j9jrK6X7uVNSfB508lm2l8l8tfeY6Tg44HtjFsZYEKb6jQxI6E/kuDCzlcTrpn
f+FB+RylW0ji6tj5BElbUvbBvXd1xOgKJO0w8LWIzHnxQpmn3TNZGnjyviPVxW9SgUPbWRsaIv9r
DDVCdztmSBk74NxPnrefTbQH8eQ984ZueTYlYvepE8E7Iy2YPuQv7U1M+/tpFDVWjd3Xfd9CbvGL
3dAKrcKPn1G5ZPTrMeqmqkimsSmgW2Yjhm2TX2YcwxFXPGVKhfwzaIUHSx/c0BTVh56JuLbQO2XH
HCqEURI8wzcwA7nsQcNA0DlxPcn4kyH0f4cXKgds6llZtMXBT7muljHmudDIjbjzg1IW6M9JLLWb
By7aJ1s03t05gPNy9c4qXZcUL2k2XaYT8Dg7apt6QwsEa0owijiKqAk7a6ykFWTMyDf4Daa5bsIB
gou4XCdah4jlzRyX98/fg2wQusXwBfj4GFq7VyRsTis97Sa7nixSDZz0jemaOyWG25HMdJGQz9Dg
nJtoaiQilE8s7a04TgICdNTrfSINS+1AaSl+5WHkME9s+te7GvGzb0hh21bEpXmrmoLO5OcrYbiS
p2LdQ6TtGDMGtRtnlHVtrZC2+hWnNPpScFVBS9FtN63WQZpD2Jd91aAYhnrAnwLiQBC4NCUFQJi4
zkcsFXvc30vcSpj4v9vhHJeKmzD/k2wlHY6JYLgEDHd4SEJjLitu/i8a1+nxnxmfgocJ2FGGEEeT
iyiRU9MC+g97VCasM53BmnsgIfMBz1kavGvmRfZ+BrXvYfjhPxPzgMML9eCpf4QUpzgJr0bSMJ7V
JjaZfJKtFmcTqbJf3abN6YgxUFEuT7zFVbK+Kt2jZUeVFrne/OW/gLrcgjKivFQz75Keib8c0vyy
Q/Vc5Dtawy7CWl70nyYGhlB+8D16lgcgCRQGiJO38LS9+hhMhXw0G/JmxQEu1Oxu3vyZpV0cPQY7
kFAATnovZa5J0ThWxWetc9efGB7j2HzUttkVAtMHgzWfKsgtVnfLQHddYqpqaDkFpvZeyujMXT+i
8q89Ec8rdr17dx/nbzke2T/wM+/0vtNRxD9a670bG7aGHUhXTCZS6IHMR9wBjFKQ177OTnAb07YU
TWn3nwJZUufy3iIqvyLHt6L9w31VOLtPrUmEsFHf1JlcQ+GH9U6CgtWWc+0XNb6g8rL9n3FXH8wU
pF7YMqiPbqPb3evi70eWFrlP/I0k+vNbsAnmoAKgM7F2KEsPi2UZIDliGeDuE0c0AvIeQwlViYQF
cEPML/+mB6hKiNeAyl3rj7yTZIHx4MKelv+77M58BLLK59xmQcFBrpwlhdiuhhuzVFAdj8cqTGBe
+JfHi9HOLtuigxIxj6vY6BgQ2BnR05oSAdrwcVsi7jdUXF64kN+TU7r1xTg+LMTzYl+4pSZziZuC
aRJBZosWq5ucvpqeSiwzNB7n0rEz5v+bh1I3h8ykZJJ3BtCBq/9nAfIstYDbbY/BD6yGMTuxmScn
i1IOliTAOG7GUzb7FMGCwBc8gDNLoii63q82uibEgFRe85Vkseeq0a4jd2CEcV6hxyfoLEU86cFX
+p1CM76fg1ged6SiXf9fXcCryu33NICybeI6QCl5AtV7V85e5nE1peto3B+bc4yeh3fPRnwQBWOQ
LFuUsNEirI/0L89u9UDI8aowE55PqUibZbRjLjwqreKl1PmCKJ7jSHJVLkY8APXvraYqP9mxZtyK
oVEhtCEAajfiTKs/DH0HHcryhZNC3mn6wV3dFRY5Pb8CoZlH/hgFlzhAmeRAq1EA1yYyXVVbdqUH
LBBX7VzrOI4YintBDwf/ONxntqntL9eqonkTsDVSzCdOBY0jodxETHWFmRHTL3B5gbY6m4jcHZPQ
X45rtAY8UWK4xY/F3r5SDdz42vYyTKK85QfkTGhiVPcXr423EwKlqU77rzhG+37iPy1t1rlumfOr
tCSNmPqOGPtVLnwfi+8y4In9y0UGrY/tWhUp7ToNCK02Hcnq0Scu0hvjqcrFN703zVJ6IHoQAF9R
WLMQpA98mDvW1inAX5DfcS2Cew/xV+nSQ4BIHuK+r1oUP4EEGRbDH693Ykp1cfK4OLHN3fFEpJ/w
HOi1rXc1I7ZbSq9P6vjiy5Zy6FyJ34TY9mBpRYM/+zgCgPcKj9cf6I2QgOe7ZilPBCARQt1w8bB3
e5W2M9II1HscQhdr4CzZtS/aIn3g4T/i9RTAC26wJdOO+SEL2ktIwxFJ1kS+qk8If7B5PUcTWaRd
l9I/JK9CyRV89aM9wOosh5FGD/0ocW5LhG7hDvkC4fRT8eJOtclCpJvcg8jaqXzGR9vqnpAhyNIs
bNU9G4JSLMenRNhQ5WtbnWsI9PSpkgKTsbufZCxV2e4kmng3EWYZ9FjHmCZ2f8vSJxXL76RIb/G9
ZKofBUuSzxNNvqTz+SLzFAKkRGUB3dRrsnIN/xxWh0yo4TzSZeAfJdCD2A9G4vW0t42xgHHZMKK/
irj63b8VvrZynXkZBZp/pffEtLZijdX0r0Gjdt/pMaAIiWZNOkD4HmgmOscQYteNVJ5mzQK69n57
nRFUcDwwfdN4djdLLi+sBMRhdAwpiihAH8fJyAwODcD5Pvlme60m+sSlN5ZMbuEHQaVDDUKTCbkr
sNIvWJsx3PFcU8LvUcK/IleRZd5Z2oYAXUkKj+0sbZue0QjH4lrEqWqtiUK1fI8Vh9MRbkSC2p0w
zeujztYKlFLNoXAIkusqeXGr88cqsH0SQlZlj8u/NIP2jdStaHVCbq3kDn034HPRF8XMMgZb+L+L
IDhdzkEaDX0Q8knBbghZEN/lVUuePW6Q/LVsP/slDM6hujQOpK9mN2gg5U+Hb+m2KGq0rUIXSoXa
QCwcT4JP4VjVpSgBdzPTnoOuHAI48hlUXFh+dgT3XPCtxKnVkzUfMiWrzYlRmHN15fPgU9VzutRa
4xN+umuvmH9snSyfC/8TK5Ijppr9d0fT0KnwAP3+Wkg8uv9kojVaEfvPrTC+EauwGJ/7HPunbAkZ
QHxab169BKBGIZeqNf/ZBrEvJVJkLhuO7D/EZe+Ev94cQP8f5/JzOiDffyroz1f2yUXG81+P6SMK
WDcXlKt3/bZJ9SeMkKzK2MgHT+jU+KyJUp4zEK0UZhx5kjxwchrOa+7E1S/CHlY6NA8eZn4p294V
YrcaziZubLw9Asv1I+E2tJ7s1FqvbdOd1Ln7NS2vgLz9RR0LTLOHgsELObfhOCsGZa7v4si04H3c
wg5O8ZBqxyzl+mk3PHRsvKxUqWJSxs3m+eHIfIx55Y6xUFKNrmVPTlZNLEna7HebzmoIx3M0BCMZ
j3f9ZXwFUUQDgR73x0F2I2OjbcHll1ajmPq4exbDRjyyskgwalK3I5pX3n7TRjQKK9VXY/ie8r3i
1dnmS6a3P3+A6MyxbGWEg+dAGWMFtr++fEawl6jZTh+W+GT73KXX6G8rbCKcruwgPS8Idw1TUbzY
Si8+JhlonSrob8TjqsUfSGu1IEA6C0GmqrxiVfdRX/catVD4HbslgIMyk3mNi7UT92xuo7HtBQJV
+FXj96Xln4FBPYYsQ5VYUnftPbVFcZ5cgFEWDmzdK5qr8bBAY+d70920vhzm4TItdGATutDCPbAr
UF+2gpD8IzZB12Hlwp0LPr7diL+FVAGCNEHxhmcEgOUOFcCoaYnY88qXz3uxbriq/c/WiXfN/AtK
IQAqmbJlH9EV3ObEiBnIzEIYIis6gmDrjj75oCvaeM0tghwCXzDRiRE/5ES90Dc7OMCJ3lGqyvl9
xL3VNhWGhjIcr4nUB3u88evssXoPvJZlRaw5RWranB40GjvBe9P5YNmykIb+pSb6QBe3PxW00pfV
1OwSpJCN7yhzvNDhQQznRg+VKgRXnXF/DL0KSEqvrtcatTwi6qCJT9yuc/jMCopjh4qvImau5Ms0
XkOOeMFl8PwQAI+t4CfDaDErJIwKnq5ce2FlZAF0LcZVG4tl5RkpKy0S2r68iIoQ3umVMJ2vLHvZ
AR471y3LWQ2170F4lm8OMuk7s9P3bet/MQ0DpLD0vzefSIjA70zlTcy+67xJAp/1RpEZAHTXub0O
ARUVZnIsMtJvK2Ybz/qZ4s4kpMRdY0S/UneF9OlQYvxhHHxRNd3YBMSGNnHdYFuSNFcHVPO8BGL3
XjlJtOsatQrC8LG3VSOej/lqM8L2hOfmB8O7stHi2Sauw3HSaNOxbNqPa/KWYmFU58tuRNJjrPgC
M3oKNPK6el3gaBEPAH2IRwqDpH8F/v0TovTofhNfWcis/NY/5s9OvcXdTWfaJtCqT8c0bPyzHNql
mVYzGe8MsRZUobYUxHs8GZQzwvlwAVNBDJi8Rhl0k5gkUz8lJL5iPVaDv05uuZoF4azRUkvFdY8A
1egTgWMMbX+lNqHTHJcZwOdwwY1RgSGe7mMjeWeCpKSFhhkwed5y5pAg8p0inrd/SgKa2UTcxVoq
9xchm1Ff4N+c4VEiEQK1Tb/9CCs2zpB88VFJWLcQby5nzVX4n8Nurz5dYiK7GFBj7kwi2WxqNvpx
gvufBChFyE0nVdXCgi+tallb7CfQRWYtSPB333N9o/6ECafpoI5/PLHbqSMG0JRfV+oDVUJV55pF
+kjZRJ+JM8fi/eMQBjFXU8L2W4bgFZ6R0x8hrPEzjjjUYihyHDccAbSf8ctQ2kRJrt8Lg+QYuqI4
Xgbj7xMEkN0lvTSfHiq0ClfYAuh7mwp6mx3LFAICRAp6cOkeY5XHSE8vHOsqmX1YnzVzGOdAE7LI
729JY/x7UNHOMk6/Y8Y5gMGVXnSAHTsbxa/D6LmzPx+8VHgoXkvpbGMVDhpxlmJ+/Nt6SrFKAhBd
7Qyk97pV9r1AqkCwlz7IUFROuuNrbrKteFFLein7R3vsKxMdeQkeuGjnYZXFJVdB+fpJydc8pFLS
CqTuIWOv3V+myq6wnokQRsmibYOFbhb6THIztUu1F+pXc+mnfBNXZXEGPNoRgPvOZUEpIJQr/gW0
6hj724q41vxpVVd8iV+7+Z5nsTPaVd8V3w/MEO56zP/hp3UHEOCpRo2/y8tShzHRgbMk0PkfKzpU
nBk3Fmb7ENVnuVNG3Lt9eG/FG99y6nq+QAwYD8cUs6/zerb4bhXnF5C7DcZ8p1KQ1yC+KGaLm3Nu
R4Ngf+vfmh6+HKeXUhE+Y+3Xa53kY0j8MQkAL45H9h/FChI6eXzhee/D58yrEdxnxG+cDp2gadCv
W1K64VhuNwJn62qc/V265gBjiT55iDRDSt32lEDRSuVHuyX4KVdOvD4gs34omukNv2OVPLwc1CXi
nrkcMHqykTzIvB1nT9VPrQKsTLQfm0OylqRinH/0tt+7nWXexqK/pmI+LebMPRzhf3oe1bhq4hAI
VUxFhY7prDRIpmUblGVnnGpuUl63B0sWG9pb/jRdajCxMwyXic1v0L7JI4dF/sQKaJDOzj7OPVXZ
0xqai8ai46OkCCZwkDTRt63q0AnkKyWokK6yUTDC0laEZYHgODEVZaY8DO0mCfVI8PuQjEYX03/8
eHZfsEDj6j8BtVmw2FUTNeYMypEVVBXuKKZT4bzB0ygaD2FVyZUp8tqRQIYdrAbR9l5cQL33ysF4
NsZ6Pfcrs2BWhjTYepp3kB+YOB+y6moxKNgGznhPjy2JZKm230W7hpzXGAbbUlEcUzwRC1CwHlm4
ySvGj4y5zCoQWusHMoD7wNrqN8eg5/idssc10F5W4Hh50DWlATRz+3wn/9kzlvELRbbFIYTBEAFd
7Vb7n9TaWiimNxBNuwdhsTDp0xrxjOR7sC578DUoBsJR04etvkPbXFPQhpWFWYLpPPQ1GiIdkisc
9RIVz6wQ0vJ934JqKRNlbm+Mi5zGkXmMl/kk7oFRjyshbMya0/qyVT+cRyhJJ9B2wIivENDwynKE
lgGfmvdX4QGkt7OL2MoYIBOMKm93KNpCSw1jQCrIeHSf1RCPERn7jd0SED8ickAu49mCCJstBCOA
VHZC7OTn3qR+3Fg/3FWnarMsGs/GxcnFQT0Uy5rUHUpGxM8TWRVmR/EM0kW8uG5dbryGbKoY8fdK
Z8iqn5483IDWBB9oxuJkIb0HEKKrg5JBFLJb/U1S/6Zuc81CIUWQ+KXgkGQcive3Jug2dmhj2Nfb
xda9XC7OrnLZFS1c9qRNgP1mO1j36yPGkmiPyoT5d4CLezCz6ZOejZ/GytZlttSdZ2dtqg+MS9PT
M2mZGLTEoH+GP8/rsgbjSfiOMUcE769p4umOGI6R80JjljY82c5vfGp6Qd/dzA0B66p2ngMo3ooQ
7WCfZkDcRRuoR/d2sFwCoRo02rLJ9+nc5SA/Yv04Eu6SuMvRFRBnLD5h5tmR7A8XSIU+2cM02deH
v8N8KpMU71eBA+le6e4nFd+u7/otMekYoZKKYpogx0mEKo5hHqCFzerckBzhxnMtLdwi0/MMWKgm
au9DxoSwLiRJg8nRPPcg294itCf6Wkuct+qgWAq6I/8uVbmf5DES6SdsRK2zQ1n8JxesVh5eDK13
fRdkPgVU/UrpEJWIvToP9H+yHXmqSEpGTKT2xTZApMcsh8854cb0pr+M5ldO7PLYDJ77RfjZuAUV
uMCWECJGWxZAPGBHliKferizwNd5/OwpAEMUqAIXfb6WHBq+PijmF7Op+pU1cEnmTN+JhfsmuopJ
pNDQbl6mr3QPfN8lGeuK/6AgByyz7FYxW0MqIfr0OpMZppiX0XB4o3b4PZgYaWgV32qETHeOwk8u
pVh3BqylMzwCuhRRQJ4I58fW5lUmFNHhv/7n68MSZDufJTSJUdSDfEwTVGUDMWlmXY/oQQUPy2Xw
KjhLX341+QXBKn5Z+TaSMjivYPKO6wxMC2bGVXJtdQtTUQ1Gu/nxXI/TbwB3AJW1ctJ8BofBDWjd
gySwdJoY53WfD2Pnh4jPGrB7CDmPejDdbHtXaaPN0ANBOVQct4ujwKUZjlykJVeR2LOxblwq4eJD
zp8FnxtxWVPMU66Ur8B2pYDbrDdzdUZs9oaIVISz0hCURPUmJ8mi0ZzpE1F3DJ6IgQ2FVq/nGqsT
uFNltGipxSAyE1h25cBADMkDlAXPduDzPAd5Y/tdIabmHHgQVyArD4cwmxLpBmJlKvl604ls0fVf
026ersJ4XrIJAVX/KzEcD4BH/Bnp5xrw6ONA9DXAbwGAdZJtlNgzst4VqDnuV0FYnf9LFdBBtblv
oJ4m+fQDEtMe/78VU7oTgZCBSXSujfo0yFhhLpuwkqXhKSzepUQZ7M4k+Xk8lgVSbyf+8C0vKs+R
fnfGs46QffZQhaWahQwdqS/bEaxE1mRx0Idont1szrWMxmibypE6Lewsiv4gV6MuN5c6/S/rafBT
Y7GhNwK+m/Kwq0ZIrAVPRGYGp+cwQ8xYoAc+fmxmcOHe6FhVeGe/PHYwVuxWPYxB5WKHE13OwuH6
3sQTd87xOtVLnETGMhX3Tlg2/RP6zUf2K8WpUonRkuunr8w85R2rUmnczUNoEYnRHLZNh0ZoXL4j
n9FOSjBzhuSKcIttYTNLml02C8sGdD64ssnOhXeL/Y72aNnzyKk7x80OlARdT4IO62lJavn+T7PF
j06OSKeZSx/0mii77BX+yIJmJPeAQ0fyWzMgGJBMNAT0jQuc3clDKlyRgGgAoFWy4eWcfFRPpEGz
HlNRm4qBV9dJKjoxljo6prOWFlmBjywLcmuUF3CoVQ43BxsbRylZkuFa+65Yp5D3nFfinrf8PnOh
BZhrSQZSHD/YCoLW3qMBJU+/OiW/bV5zLeB5Q4w+t2UxpXw+4S7llDpNGOpMBQh3ehcGJD3Du7io
zo/z7EMMnkpyzl00nHSxipc3PV57ujPnOIvvXv2XQ1+BcvVYyoj06r9I0HNgGLVfKyNoy0J+cK2H
SAR3+QmTiZd5DnE5Zd7CZIgE5racChMbwwjRLlm0r7woUqIMHkDKIppaq/mM6ZmD7BbTEjTIxmhE
UtmO2TJE07EfMFwjikbFlHMSaBoHRyqXHT0kCqxzYddv0NhQihxMrKUMVz5m+AU+glGIugd5Oj/F
EBdyd71FWz2306d6lZc6kwJP+SLPfyWOJqGsTmhBXQ/p1QWqR44M0uaSTPBgAimqIoNItsyaTjQ4
EzaLZ4tu0oO3kUxMqg8SE67YihPghGIYk0Z8WEH1gOmyzbQhvVk/FkkizLo6qVI67kqV053ekXvX
moFL2XA/ten+/6ZOngEn26NeCoxCOznoJYCzFgJAY7LM9sKAwwHLEJVARetjGbRpicfrVEm0vT3W
/SZ6ao8yhdB1phucIGha1lgZqAAxx1RQpJ2HaBLizXIig1cMejfBjF7ZS5naY0p718Pvpqvif59+
sNvKa0x770/q0XadD61qwGkMk49CJbIaIlVL3H9nGz7fOpBx7xDqXLv+HR7U/yfXprfpcjszQ9gh
hpLPTugMsztDKvAo0MsLKZDpcrJXWfJlk/nBpIRxDB3xT9LGt5p9aAtJmupJ4WT3DDYY/eZiyOH9
RIK9RhTBkkZS4d6D41u3oU5cXHuzlCNEVWqGMGqx28nv3Cz83oW9TZAxXpY9wqA+aMm4RisZD2h2
AEPBeTe6QFLYZmA1yBP2H39eZf5knKAJbcRHfaIIEJEhgmtdZzR+YS3npaVp7f2h6ow9H6qTCh8X
ixZe/MQb9LjhQTbT0vwtSN5f84qh2WGbrZxgxCz1TYM1RruKiXXwdk9vtjiMjtZ0FU8qcQmIrMBV
fzo5ZzlPWxbb8sE1I22AP38qghDH7oXYs8+mZM08v/UHbwb/HvZnVTB4YDnvDXDklvaNcKWabY+8
pXDweANA/2Dx0Nsr5rBLTOxYeSZVyj/FrkJXgBLaigz0Q2g1oOKZ/Y+ZBMZO52hX9m3FeCXtDhDu
bNl8BE263X2IcE9sUlcdc8BJhxEdizG7TooOhjEKj+LnpblBTXoCHQm19wLtfYelntTadEUVJHnk
Qt3//G8KuYlKK0dcT8PGDb/kwltMQoK0zXQk1Zyvnz+asIh+B+pqXrivgCHMiGdx3QEex1RIBl6R
CeIO/BgjwWvIGPljRhE+UyphAqA3BpCahnidKlM6PoPX6HZr4ejee+Wu6WkstPRB/tTq1nAW07P1
1fJ7BboD9ctYbbqN6Y6w0gBny2sMfntHJ78CkiIcU7X0XAzS1P9WL4kFxKEr6YoJCfaKHL9U7OGu
/SoJa86fIi7huW6CvyFeIwUgiuleHq8qO+WsD9YwUlce2oaPSjkL+JQGxCJ42ZSAlRCECFmhKzVX
DzmdkKKeP12P3CPmkPKX8m6N/2iXph+1G5BgU4jPWreraKdPvvedXk5o1ugc2E6P3QPupXgWZx0X
muXxPIcTQdGBsU84TBvPgh+EfaZr5zzbImDfBaL5WcZ9U/lOyUJYmyX2KEHWWpxlZMcsUz2oNxvt
/G+wwqv2MnbTQnjMt1TS7eRy6UxOd0z3NjebdkgdFUaP8vJLDOdJxZA2Zuv0A2Wu4XR19j8tqHcP
ZfQi8CJl/wacVtZBtXehopYH7WouV6+Unip7HcoiHKPW8JRSogF4NH07caKr4YmoxydccJnqNVGt
qzsxCpQ4vNhfmAWjuc/gEZJ+wFogtdDa6H2TjXVAn5Lu65TLvyImRedXbKZaR9lUqWqw4y+zdWc4
1Kgx3K285WNkWIJd/TVYbWi02z1Ss4B/UBVmhbC8jT6RLnnbkwUDw51x8P0mdhHO+A4XoRr7g13s
Wix9HehWf4SshxouITNcRfrjQxsIwkgjGf/kbPsXFTBcr1Gw5zL4rXmg5iIJNtGd6/23NsjNKPzh
CxQbcvZkjQuTFUOszBov92WA9YScC8sD8pNjsDeLpnPispbDGA0dsecdpNhymSelivOtO2LDz3av
0j949TCQwq0CqmXKeA5Q1DHbuMkcm3UrDFVvKsuAkOzaWdfc0Xczy+HzUfl5WX+r7zPPlH/rNZIR
cmfrorXdC5WSj6ExpZwsggKY+HE2MqW5fe6kO1eUlRvkxFmvW8H3Lj4JK7yL4t/NKyU3x7GU0PCo
3qhlkzyYv0/gYm30C33LxWJyiVHeNqLGccKOw+nBsmymCyx/fXhJHe/S55nogwpKo3VwG2yjO2KZ
EMpkfKb0zmY70jv6+gJ/3XMUlGiRczX6Yl0HPfLe9MEKRdqiQU4t7n//cas58OhQsPrHcc5/AS6J
B6peNtsUoJm7oD/H+gkX56g9xFNWX449QvRS6R7xWZZ4wy8HQzznTBOFHEiYnMSApRwBBDFJnvbZ
2vDP3D29PV48Mlvfe8LogO3+LhZGgKN6rilXIdOJF1qu0hIz3g90tbQ6+buRhNdaCUdgtNTXjQsg
R4ypcku8qSqN25roIWsoy59iJ6zXQNuusnUM+jA3MEkH4Y+edsgfqnRi8CpASmbvRuBc51G4SXy5
w/uLPp1DM9HTq6/q2B7rmnMeHXWabRE8fwoYVyNVeqffQjWVwGbmJxhlXeQ0EdEDEElV7TTuiwc3
6kO9OqEg2Ay4A7bOhAAfIfsgziHrYi8OVB3TOu799ASArKxDEMt5o94FHk9YFaT09m2U0H7B/fAC
JXJ8mALFAiM5wYeHHm7bw/vg5dKGyl1AYhfYx+xoj61ieDLIGRZz6QLu4oDnbbIEy0uvhsAWrsvk
X+SdcWG4NrBolX/KW/D9hTytcOwWkLdJvuKJZGz0KoJ6MSz2TE/r8L5cntZpz7DOccUfytmL2ndb
bRac5RrCKs+EXrUw+auSebZqX59mUOFRLp9GNdv7rxvTEPj2yql5NuNHzJqohLeHvhu4I+rCnkdM
Oss6LaJrcvyxgjuD4eXrW9PenACBbC6/XCt/uAkol1Yd/bDJ0uPk9sddzZ+AfzU9Zcr1MC4d3C+J
P6ARCJLNgWxPk2bHMmLtY22Zc7946IFBMbOeBVtd2atnQaeSy71LGutXZrm8o8GaEpwr5jo/tInq
2UEKt6w5yvzW48pYCHElRf+O0TFZzFSCy+FkhdlblTny9jwMlxIcTctGPyui69j/mFRhbt6Ai/b8
1YWUoW4w2Tf6h/36uMDjGfPywtkvpjpL/n+6oIofY3mUo3cv4RwHQXcTIVBHTsavjGX39N0gA1ku
Z2QF/rvbf31qvfAqI4u8XVgqyC2KobF0za8m4EcIdj673v+ybubD9MdjBaBQEeHT2nWnVWwD6IIn
QsHD9RrKNll3IjnTyhWpTRTBnkt5fNbOd9L1CBRPYQe/5RqxErrrQ8/d1hJ2QqIgo7ZXDfRuOj1M
aqFFbgbjHYCCKrLxCDQ1aeJSJ7flbsNYwr4vPZUF42BV2oTCgUA/dHMoE+25iQlMIjeG3LqH4/r5
dIIXcK7rHPJvEJ2n2h2MhcSMlRuQuDUdplL3yWCTl6H9WNLxN8KSr6jg6/L9eDapt1Zhwdr6HuWK
efAHNuvr5Ic1nY6IS4d3+oPMpd35WXh5A9Y6QiZDkGRoIlm3TWtSDzjfdCPDIs3fehVjlp7oFMN4
TGBQZgAIb2v0JVXk7K4TdmYj+EHaqr+7gtvHwhmHDW6rz0jKez6yyXAwOT9thbdlrynnIpdRf6zS
oOXDc2VXUzck3pXARerGSaQLm1mS8MHEl5oMGcNOyDNk4tHcFfzTciwjHmM/m7jLPAQ7bEmVxGgp
bs8iPiQ/ACRTC6agdRfrZAomGmz7geocFd8uPlF6a0wQTpjBOlojNlPCcrF+gDBLZMCZ5wd8UaSR
+lp9uk9nD6iNqpd6qVSmrEi2NXqBc3rXOpSww2ZNiv9A3vmwzz8oRI0ISfUxj8ro5YHQDMthwN2j
CIyd4vIUkCkXY0jOPsKMZWwuZ4VwGbfOdEMmEuXaQuIA+8hNbeiXogdBfIUEAtYsoUOHi65qTdg1
3xpgLW2BeMo3KGPOiRKkwk+u8q2ZIyK7upn0bVOLqwsm9L3q/Im04O4YQpcsK5YbTXom5nBmTzAK
4AXtN21XASyj+63/xl24nSEbbOE4XnwWysSlNHv9YkUoeh+s+WC82UXfBwydv7zIzsFRxrZuZF+G
DX97i24MtIkMOxNruX6YryH9cw0Cu6zlM7sOpmFdGd9r4A+7/gqd1UH2dUSeL3tXyqd3jMguKcIj
SM6lo4fASJFHkbi79qM8BMXQ4mNpwInaMSVP46EPfijLD8mhBTLQ3zUgVXplZsJIWIVFKFCHxf4E
Zi6ajwB6AKMjg4ExGEW6vdPa6A+CsZQINopoTn5AKtZ6bDA7PHDQ3vc6rFMm7qgwLJGYZ2l/3f4O
5hVe1JZs1wmhJDq7yHZ6K5JBqF6asTgcY4mAURlP2lgnnU1QgI4KI7ZR3otYyvrp+y6l8wuVkVZv
LlV4wAMgRWQ4F2TPbVckFd51/5hatb99TnAbsXOVADTk3ZLiB+N6zlS1PxJnloYi88LPD+IYEoKh
AQTBfxh+Im0FG3TibGoIRuIYHaRgIqY7u0cNzXTzlw0zjo1PumRMpJOWMFBiEp1cm2zmopal2vfD
p6y0GONjAeYHuax5vMQXLnH/dya8xjAK0fMOj8DVqSIbeM9y062zt+i9ACUnelp4iXdLGFUln6h2
F0UdJ8o41hh7KXluCaAg12jJ3G7QuO6vs/1hDiUGvDqX2HOdUCs4KpybZtZVDH3W2QgPB7gceqzP
WzXMYgQFd09JwaJbG0DewYiA3Qvzr2aHdNBEdYr3g7tM3uXi/ZrdoOZQXp+FK/QDAd5SDt/EgSpp
NIGJSzodzEYwRWfTshlPHBWjsFHrg55yKuhMEuWMODjlITZxAJj746NxbVDD9d293ffVds2eL9zG
fFz17ELlLWpTz3hR/aqJjUo6Yy1mTxJta0Osm3O0+NLlllZSi2Fzc8jk5bW71iXr9cIe4Qh0bbhT
igSRKoj/HDDcGYLmKxwK8WVW38EMYIFTT+VmD3F+KkVZfC/vgb5U+RKDwkekWC4Z76Z0wLS3Uy2c
ZLCWh4OxgujCcv0vyA15CsSr+KjUfO087b5R1xV/e/KTFSXVZsPWK3kiM2a4yJke3YTuTFcdTZ3G
JM166nPTNtxMT3rXTqrWgLTvyXRr7EKVKTjj/llUPRZEb9X3gIRpYKnFY4wKZB3cADwqRo3ToZ5a
lSwiqk8pQjxVbmhp/X/rRWoPtCI9ngLMBDph9m6Phz3hcj0UmGfy2xboqMeg9GEG1YIwSeAK7hEg
YoCyZ11bQlpncqQfTKtLcDf9W2u7ocLpV/8n3DUCYbvYVPeXKQT4/uR4xZcKWdajs1YdsuxdWVxJ
Xir9+KKrbf2UtR9C1bd/eV9Sp4EezLojohs34edq1oJ39KbctC/yozxDVK0dz2yVzEaZKtPZbWB9
ou9b4Z/wAJsV36Hp3Ze0L4M1tsAfM4PtpznntGKl2Is3GKlJmPBZoQAzRIUrDevHMcyUZNZuZzMj
3qgLcePcTUVuHMoHp5Y0rD75Tr0HbFzY9p0+q3UgcByU/in4mqo2WT16OQjou9JTg+s4acEtrUpS
btJseyTIOBvOlYXDrrnmWp2d/fyoqDno27VXvZV7aDASZLy7kg+d2XLDtrbcNVuXa2O4npqAuumh
BPDH2148ZLhLbL98RRSxAWC4XAB1STUCLuY3NNT6xmau9zqEG/HqygaTu6xOMUFN3kJrmm3ZlCqA
Tvy47x1LrjnvFJ1r3CcT3JRP/hyIA8NOSsbdKJk6RbhpVpDt/WazrDti3bEmQdjMzIh8YLpOqvA3
lzQwT3dVmvv6YOEQu8XR+YdNxkbjO1pooeJY++4RVAKyi37XNKReanuSMsN5p1684njHYB/4IvLd
0TGHACpJEQaWrA1tbaAP8/P0UvkAk9tg+OK+XGbYwjk65xUBltRBNRCAL9Z8FQlp0NWaz4MABtCj
jyb6V2/0JnpvDA4nJzckkZlRKoisTmCIQOv5na4A4ppT+8RYb53t4+fmElXJZvsaujE+LtqWBWuT
T0fuOWbJ06N+DlDQFB0fjs6UGoFZP/ZfwSPHjK8zTJcFfPcHbBil3kcnUeRWotlYFbttBoapK7Ni
yUTx89fU4q4cyE0lf2Jt1ugJPlcakdGOYE90c+snCf4xGQ4=
`pragma protect end_protected

