`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
j8rghYExxugJ3wDse0b6EaeS2mTwYZtMOIUthb7h89zRBHObVhsPjtsIS2kXljjtVIIiBpoPqIqB
qlGHzxD/L9J8r/XS63Pi0a1MtYo85k0nQjj+3YfVtHKnfGmPpkCaxf8Y9cAcP8TgfPvrvJIg5Q6k
3BF998YyMyIDuhe4FH2kRB2c1O5C9lpQyaLUBZ6p2GwwXyiu69TUwKDq0VdxR6fxKwu6wUZLa17I
UCnZBrDMTSHc7TgAkt5OeV9wqbdKV/azUBR4tjoUV89gu5q0w48Wj/IoIsPbAN/I2X5S3I67kuCn
V+50tmhfbG6KYo0og1Q8jRsi+VZDQQDGn2mnQw==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
ZBwiJamtE7re6E9MnO1PlBeGJ7JPNGmISlzREdFr3quxNCzbEUesc6dBx7MedSJbgWRk6gOGxFgx
WmSFteToDQ9f+7nZ5gKRsxwIH+3WcEzZPmIHsCBbqqodZpJajB8pVCDPm9SO/jiKFnt+hoXDGKen
8GVe1CaBZHpK6maLwZwC3F8iMHMX2HkJZp0rWtLeurwrawKFKvymJdqMuWNhAIJoCzCp4QhycqcQ
r85bVmQV+ljB0wT+l7O3Ss2JE6TuPzkUZKtkoQf8d9lIX4PY+3foDRjt6KXY2LXAbLd9hu0vKhT8
iJP4q6sCXlqizNrT2rkH+7ui4qOkblwtpk+fNwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
oDYcyl2/YKukWyxMJFUZ8FRFSOXBGXEPT55GZEM5ZlbPEQgW9irnDYeBPH3R2LAdbjT5mqfIMoAv
KGCoadUAnA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A+alMHaI+s9d9NcU6z/cZbVAee+v5L4yA1vdrOFPjn4o+za4W7WoNtR1c14cD0WtJBLQrA0qWt8Q
hmqiZLa7NhQF2oOC08bimSSoyV1rRLohqm52VQg//e/zb/zVzNKz+pOjYS7uhD1IKfW6KfM6UgBM
jGI2dTWXTrkBYCAIQtJllO7RtkcQ2JTtcd+hAAGGKG+s5Xgf35Oib6RrCoxuHjPE4KxiApSyanrF
c7lEAVxT5GrGy5GUYxd4oHLJ1n98QJtk/mBs9HwmPXLvJRM8LZFqPBSpdd9X4rUGw2+CbAVSS3pX
T3y9nSj1XZWprBX5AOLGbM0cA2U7SO/AZKdgig==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rYLjXxvKZdOcP3XdyBK2gfkjCF1E95ZL+PCvtzjx6xHOKpdHE5hkWL3W5fDChkHNnynz/HV8x13I
hXbqd1zzktF1uivxeMrbFG9WsriFBcYYNYFAS4ElNtMsuD2aMx383FsXPpQWbPm2+gobIBUpBZH/
/x2Wi/0YrfyG5o5yPlfuU6W10rUhXaGu3cHiRnrgW6L72oG2zh40QHpvUcJEa94koL6e6uUvmeFn
a1p3dDxcBJpGeBc9g9b+80Y52IBd2ZjgdV0DS2EfJBzuRvWZF1X1Ah9VegJCLPGbKIesPLLXAuk0
ix7bSW+8MgwjQcbo/Nn7yc2o9zB91MvZB38BHA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DTT6NnjX2RTAInegjUQeaqobCtQZ2NqwM7cxz3MHjDmTfHxGaIGWJTZczk3qQBzvhAnDZN1oBFkF
Kjt9nt/n1ySQuU6f8Ew1FQp0AO1Var5HJt+N7VetFqk/Awg371osGFXio2fH00OjMglAhKFRkeFx
Z69wJBcStLYEMry/RhU=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U2d3pmM+us5NuHDrLVSsgLBalxhOBdJQL9WpyDrhUHmvvR7it4kl2PQpd7hyN7+jO2SdY93njBvY
H3vGTzYZDIbemd3mcfF89kVCQKIhdjzn2blSdZ/xQx1HZOfFbZUFddhBw3fE9OCRm/oP2+Zmienm
G26Ncf3s+wcMxpF1gS/VE9466B6OHwZWkMYWXifG/YMRbD69qpg+1KQpqcUKeP3tgodPT0i8CX3g
o713I3nvCHVwx3m1og5xi5XBu5ndjN4X2cnrRuMzoyKaMUAWCnDM9wm4ezOHU8bOB7iVea6c+JXI
XQYJSuAW8koZjJ44yzCKvIayqoGgiqhzPlwJlQ==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SNRNeVS92XOcf0USDgWQL1W+aRpY8/B2NLztV3MHzYM58sYNrLbyDl3FKC2vTteeMHsSRrcuwZr+
PsTb28NT55PwGWzvSz2bvld5N6d2Jor982/nVa+0dsLr8M4YJ5sXWDKdK9u7imSkCwlj8f6ENS/p
7Ua7WEnheSTSSQnu4s6L8429Bz6M3JgVr0V9VBob2OE/VB/DIWuOnl5RIYPk/Evl7O7JvjUu62AO
PlpDaL1YKbFAPLPS9mxTNbHUScABMVBTtuUdowrq7iMIFIpndKFgR74vpLuTuVMBdjZgZps/TnjN
R3BRGGuD4Eiitu2IvcKG++qB34zLt0cXA2baZA==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
H+ifCezats9cXTzUnjFatunXay0ijOWJD5pGgZDKSbyZY/mjpGPFI/Y5mvBLj3GsIi55X8wy/OxN
4J3VtB8EnbcbkuoyRxI0oHYFq3J1/7EvrN3XjnjSIkHTNZqcPeQAdcnrenFGCGBGrUuW67VzZd6b
dxvyvTe6C1iT7I1FWKA=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
EEohfe8vApfjeu5136jQxQFFJV9IxLuKJYf5RpgFFSxot1GY9sQ3IbVpLPuosw5De7+Gp64kGN6Y
a2Hs/F1rEe2YiGZMJiiqOfH1Ce9DbTrbvEnMxFwLQNhf0Wm5DDGCMkwKzmDNYj6TR8T5UI4Rp9qE
fIxe4Zr9hPCU+3lzY5BWymYA4mLQ6q0SREayeO1c52cVdpraLoa12eUo+8EDVlyhCqdM6ehmHeir
yP9nmZFDubiSXOBX5WJGVQ3X3DzubvUm5KQknCmzo4hkqO3dW5uWOJjYDZdFvPfeKwrUmlAkEkDs
c71NGYLgttm2CTbtWvuhgbTKB2aXOXnuDe4F6g==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71312)
`pragma protect data_block
6dWgl7VbtdcBoc9kgbu4Y2cE0CizTLe6mtNIq5vORpW6sd8FeFZLIL0/2UBX6Gb0b6T7n2n70lev
ovuEnsg26vVW3GJGCgaL+bHI1srOx1tTAfkYG/2CtzZaoUvexvltKqoYlzA60B2JFx9/VmAWRIiQ
ANwOwaI7YJXLN9a3WfPeGj93yDgaBChrzfeS9wkUfNJ/d50G6bbYv97VHe3teqOm8ciiuc3aZUV0
0bq9eyaClPudZRTuAuAqAXZ+Nf1OVj3nONw/HVxqbZ+PvD0E8g9bWsjYVt+ffPGHR6jKbPy212vH
1RNRuFgY/SUkhNmW0jAE4mmplTxTwu925dv7TuPwbYTmm7Vc6N93+FSVKyEVxcLx84lOEN90kHC6
ERCOSRb3l+rN5d6Feor5DgzU+4M3ZMrWhTo97xWXLVWAPU8M+/VNWwC3xcMQDG1SarvDI65J6+xC
IHjmULK2VueDprtEcugr8p+sz0w5aCO4mTTSrq82+58YQ0p1Utgc3i8OLx6pOmotGEwKNmO8IS8w
+ULT0BhSUYNDcPaDTxSpgs835bWTKiQDowq1i8qwDWnt6Ha0bG5B4tPmh3+NMhnmL/99TcKTzUTj
bcjQV5Pj8WdXrL1u4tRNhXL6gEZW0eXUTmN/vbvNZXOvpPC598puQ7X5Cn2PISdHBSp7tLBQCyxl
WgD2GYi192svZpILxEVvpQQLqWciszYWNrN6z7OWxqJSrn2Ih6gVawgGNIr7Rtwt7nX2XEvXdSgW
5gXBn6ZgQ5THtsa/tCkHGDv311NmxkRPUXuDK3u7V2zXPZyvqBm3kKHFXJJ6ipWigEvCO2YF9PRY
kYQeZtStlI41er7yRzoBdxv8Jaf+vDyIpRmBPz9fszAZZOPYuAXwBdiIi2iqi3c5HOX76UitApkK
vp3+lHutHj8iRXfBCFyl44vBAc3ZQX5XnDs9slKKYYiFs8h2wuOENxGOaEMPMzfaoHqqtrHwCLEo
wrtsS9iEST/B2DK9TwgljWLN6OsthmQbO1U+7ANqDaKgOWTPJyjvsO8yRBD/2vNUgoDyNJy16a7K
tmRRAJxoogEEtEibgNDmsqZexFl1S70SL8VDf1A1NIzxE59zWMm+zxu02HfmxFjeGBNjkoEC4pCA
J//eFa8PIpKfijFx6aAkAAyYYmF7+EvYSBLHFzMKFItJXLANcYat/+QZNRU3Qjt0gFej4tYwjdkI
Eo7UVqLuVNf5B0Q5ejHU+e+wh/htoyN1LdfPhdaEMdcQ5pOpgBmsVYWoNpe+7/OV5H/T/VSnAX9c
L/aJK6w/9B4OD9tZsjJ1swJG/JPzmRlhsbsFFtnpdYGce4NnTUyRS4rC6WKvVkmlObqF1HE6pKGr
hdFLNOcnuNghUmckU/Sk/KWMAEnTdNQcNdhnZLml0oqwHyS6Qk6uRXSrAJ6jXhsd2XgzxBO7e3EC
kaIfNGYSsY85RmxSfMZiANf2lAryiKJH8zKoxf1wAMZ36wKrAoLvPoltqSPfTj3OJV14hZkH1t2Y
hNnvTxcYu84+H7wME+5Npj9tXphP2Jim9Qpu59Ikm1qiz/iTFi/dGCheOevnpsCnU/KnmVOZqcjB
keOxIPYBvBL+UBGvviMfHL45PhBDX1AztcdvQqDrY3PxWHBpHfrXlUHAB+Nj4HiSTZf9f/k4Kc67
YHKHXhNelmlzCBN/nSIV72g5KVIeiUqsorR8cLFST+FfIqoXdiLPeQOuIPYODnSl1lJemKW2Kysh
EgGQZlzQgUS87xG1jS9z2j0mSY/kVSsLymjH5WKvdK0r8Os8OPk0GtaPfvCx0ovoHURD/xdUSzNR
FLOsPo0oxQKlljdabaNYR6McKO16V0S4stgW3F3gg4KdqdsuLEBAIavTFMX4mJfrd2q+ldPCVDQK
3v7esK3Yw/dkaRhOMAsZtOMhmx1ycwdoggbfCVdFSs5uWhdLhvg7PacVr4klzu8X73d08gIxhdiT
wKPOHCXpnWD5qxHLzHfoBQq3YNQAUs+nNo5g8derFH0dlJe+VcwrZWVwISxdjDJ17x1XwZJA1AgN
a2zcxcV2gWwjioARyb4M7OyF5CLWu63SKaH4TFvgfMAiSh7nNJLgrofryBSlLna0RFNvrwC5RFQ1
F01MpTZvgypVa5FMMpoXzNQe9yJPRy/0AkoKMnPVnEnoPUrFRHnUlGayb0TMWWVmkfX4oynov+GT
PezPjP2Em96dO/1z9utcB4O3Q7NHYWOwaLsqWKwQI5cKCuCF2xvuVVxmWczlU6sPs0irpPK2vaA4
Pk2gAZEA759UEU+lRtk20PRCalHE3bjzdiZwXEYW5PA1jlIo60NVYwj2iAXop+ZaLlbuHNQE4zn8
uVUE86BZTMaaZ5fRrLO3pbvOJWrczvr6cDaSWAgRRB0JzOxGyWIw1Wsu54XfuG52Nkg+odywbAMm
vxO5ndg8G7yrDJbiyOBTy7VGaYgHiaEZIBCR6U+jY+UlnauxeAoc1HXsz8vAejZVVr/23DoXe0bc
a1KyYL4VHwa0QsxVoY9jrnOdMUcotxOjpONMPpmSfIpxPX9EwA/5YFIK3sZjMJj8CLOGvD8+vqXj
kw0qk9lh6BN3K77GgN1CKDwgtvDaqJR3LbjMbRdf+oin7d2CoZj8vsR/DmDanDzPairkS6mEHAeX
KhNKUFSb/TLL+pOtC9HRnaKp/B/bFcGEWL6igzF9mDxZ1AHYlHCjvblYzozmHzT5zwUnkQziSAGl
XMOGuw88uMLZPO9eUL8h3e7F+I/f3rTM4Lco9WEy0hJK3LAcvQKkHzOn+1Ja4xKXe7WRbsN7VOx8
LFVWMFHjo3bNeGdL6spktJYWEbjfKyqKYEFba1q46NqifhoYzaFkeGcqa/br2legfnJYsUxOaLbl
b46PC0r5pbbwA+yGq9B/Gi+16yLUaZ/PdZNbv2WBDBC7dA7I+m2VwevR957LSto/8mNfKjEq8jkX
ticHkhPgwi7EVasICjYbfoWLRGAJDHTOSlXGaqWeeN92CHtB4C81vJAyOV9/WYVMQkR2e4aHXjdw
CnrLVhknD52QcLTsJcHrXPlUUlL3FA3w6oAYcrHMDuDY4BRs8jE/WeGLMNHxviRMKFV3mtqOQ8LT
z9ziPalLkXgufeanZWztTv3uR8LXdzv53GmE3e8SEyWDLMSOF7gEHR+1cm80CY8WRhjURd1qL3NV
F5FnNIcHthnuOjtxd9UaEFYfLBxFSCAjyVeY7+4rRoePP7Zk35qO49zhMOIj7JZQhbKB/gNOlOkA
Ogsk81nn1VbJmHMoeLcpFmUmgVsdiepEgsveMhTsxO3ydU5DK/TTMPev7dPgyipM+suzSEzDWDuc
I3pTNeLnZDDIeuWjMQyEjtEy25VUX2aiGaWryKiGE8ww1A8zV2vqENpZZekKVnz1SKnfYQvDBB+1
9xSi9koShZ2kQoZeOlhxWys2PWux7wqybhUzpXWkqOsmL6+pfCQ9cNVpEXat+vzOzJfbjeh8K5lF
dhvefaAbRjYaI/MqDK/8IvtxhBb2lbaorBwrOZ6YeWaxAKZSoAD7dS0iuEVepE+GopWDfaZq301j
wg5qlm1+GEljCTDVlllLdXq3GkuAXyla0QWvuOqojN4Uym7bZPNRfO39fDCyOssJGl+aSGoju4Vf
PELFBOiM8rYNkqySopwA+fkeVLjmu3JtTFyIHmJKDY4Vb2coyfOnjdWBMu3Xl7kJKuemcGdBaJCG
nMwgbF1TpI7GscqdJzEsMO4E1nCDoeTck7/1PZuREpD1JI4mES76W37rXx9OjNZrpMuCSxmCe1Yo
jSZaEeejDmnhJSLIJzb/IeaNF7p7LRE/RwgB9kpgWayKkTcw4hV4wodRYIbq/jImEWzs7ZyW++GO
V1DLxdNMCcQokmL6Ujn2qpcNKgywjSjYQZKoASbmVpxrUcG4ezB3RK1LSZnC7eeOd2C79R6gR+vS
/nfinHeiESoy1sHK8/fUR+2kYhP7FgHLqsrcQoOqjwphBvRIPtPo26Ptcj0SxdQ3fAXWe7RtpXJS
cNeuhAn1YlH1fry/FHrOXZG2qDOmfXgoQKrhFdjr/eqt2dhtK5JcUH+N1CjYO33O+TP4CIYn+aJk
0LggAq2S8LVOXEkunHIQYIjrksUns8Z+LuSr8yTE4pKZ66W/LFuEGQIjZXZ/bCLeN0joNjnQO8gq
S4iQPiNlxzHz7P1iTnPU4blwmyw5Y4/RDJhUeqGYkP7YSY3WZq1SAduqzLYReRfIENhHtvzGvpuG
xuUsnKygoHUYxRCPZ3yCVPh4XWwq/eLIC9npzEtNxf004pa6DdOTmqHqi8i+pLUqyzXWr/kFHw5L
RAwni1u1i14meovrWa9nMyJi952RGEFoe0zFyNo2f8JdT3zj7Ciha2M2Oob4DIb6ZLvXoLsh82Nt
3tAagA68M5PnldAy72xVwwsOVQi3ei1j8buoJi94PWcETwF2d7d2HfYvfDE4CKuKBUs3ooaNW03G
Q+jNCcxDjqWFxRmDIbXJxuqqZnb5+N4JOojMWqedQsDqtF4VMGw9ODvQebintEO8d59JlXNGPUnO
bQGbUIk9Ni+gPwYtPSxFFO3Xe/DNjCmo8VkOuxh86ghD/RgxYkMKopg9VsmfuGJdaChBIHvXBIg+
oDhSHkMokzxoVfgHQMvqI5RAcGRs4wMKLo9Z4Y+jqPIAwrZqiSKYGskZPbBUZZNvN+g6c8jjjsum
UQ7ITrBcKED/Zj87Oa0vInAs13kxiNqkFHu7n7av1spN3LlnVn3pxPyWfVnQ6ct1l7JOgoqc+rfk
+8VEPHlz3oT0JHQul59xBy13Zli0Yf3uMEkxy/Xo2/4FzvmusIfAvNpk/cbilvavxQF4tdGU6lrA
wy34cPcn7YZExT8a4g0z+lCzhUpDbxDeghEmXYvvBjn4chgq28+fFX34m7a9J2WJtq1aaxqwgGdD
hDLRsp5SlZW7iip+4wTCW2VrjS0gMaWYllCfbbGn2sitKU79q9cYvCCHA/yq26BKVlEYoAsmJhZ+
BUs4yBjrAGftl/woUxGyJQ7lZI20NdzWTIKwXHMwXMURCXXTo8HSLbSDhBHmk/BUPtiQJkMwzhKH
oQP23eBKX1akrntAuGDJTRReiV3lWyEuRim96MrbNRqWUATB22dhuGX3QRqVL72Go3fu4hQd4WJr
Jss2XWO97b5fWTB5JS8NQO2PRhqThpRmh604RLfP+vLOVRwCGnlMKN56qIUXPNt1GQCawdRAvTTe
Lqq1kcrNManRVCXDX8o4CzrUvrU5Re5dL94BzS8Mdt6kUixjeX0CUQ2Qf4KxSEe7WUg30vCI0ugW
aSsUuGCPK7KDq3Eq1wucoPWywgKq/R4ZriPk0PBcoWpCSxA14GGkDDRLGBG3yss2Wp2DaH4cdlYX
BuCK31PuF+AM7E8kRR9bklFzjH3aoQ1fBlzKTF1I7G6nZ/lyzTodvxhW92a5t+MoTLIaAKhztb7K
KibXourjaRbSEZWRPfx1iLUHGJHjmfsNiVTw05HUbip4s9Q5C6TYYv6AD/YKEHTlk3vvO4rIwdL5
BNen1PFLqq1VU3SFtvpHji4o5l9TLkJeEaPECekub9mHGy03cqjs8mz2iD1C1cFoS2LLK5ImgO5g
ptdL8GT9oBIwtV5HyGlQiiyxiIB+X6hxocBDdm7BOnSCZDgxY9WyQiNtgOUOHSx9hbdyjnLVwLF1
Ei0ZRzSOyrki+sQdmBCiCZOFfHc5pIpmRh3YaUXA3hEU/Ft9iMzS/ie7Q90yG3pnJo7kVYUR+BKD
4eW0O2tggaXkuex95eWGCD+COf98+wy+w9uCSTK5O/lGwwWzmspPkcSpPwEnT0X9o/2DVT0VtLpv
py4+pCRIqrafGWewLRk+wX1I5He8Lkhg9UAHdCvLPtwqa/0G95ADHiDGVpy7S5wGPLvBisu1Egyk
o2XDytTArPrxNvdGJo8EseTI9yjBWzNYrreeYdf2mS0G+XL8naGR+utzx2Qaiq0ldLbpt9bPGkjL
qurSFP9tgY9dCwMfvMtm8ZlxfHF5LZjju/ykuRo4/zCW2CSm1UjQXccC04PnSF+e4bW0+6bTQR+B
LfPKva89xJ9hyQOayyRwd4TpgscVjV2MJqRv057QK0N4NW6kPR3+uPYAFruBZpDLCDGjeallVD2p
3Ie1KqzYIZzOsIiYYj4ONW0l21w9DESHESpohk9lTu8aYD7roveV2UrN2vDHhPX1QzcyJB3UxFVJ
IZysquxFqSIxGV8I8cu6Q8s7P0f/7cVSLLUCGbwIU9Z2p5GqPcmPInY9IfYgVF6XhLItaXibR4uG
BohGAnZhPYphB+0kLoIApgLS/IT+e1E69c8kwUSAeSpTSNAJR2HZgDswku+tuaY6Ltjqk7Y+Uz8C
ouZXAszzwcdf3e/ObfDNcMKkucx77ZYxBEkGaE/K6a8B/0H87bLfAAvhqaP3MT3qPx4SIbn6x/2K
Zs7XVtbPs0biCLdK9z+hzkTAgP/BqgT1scKD7hmRqzFeKcqnc26PzYapoLC2xmxM31ztFMv6roEJ
BTXEpOXx2W9oKck0Gusf5bD0+uIyu0R85ukPqSnsriXcT4myAbHGQMJu9hVhjE+2R5kbsbSfSWTY
r22NNboNz2huAR5TpcgsKKzIQ+9yDbKSUD+OWwpASshgnYRwPCBatdHejLiXTmXjYK/FyjeU7JPd
fgKYrzj180UIWRobWJuU1AVNlQL/YP0zq1vlMOkghBN/eYSvzl35e0c7V0VpArKjm0gRY1Is7ZNO
fy6jysiLIZm4ApFJQ8cxBpZw5vfJ2JdRf7eoo4HvBC89tGw9FQ3bVDI5RXO2+iqV6n+5y7N30Qul
pS3ttwawDhr3GmZKKjBMgR1THt+8sX5OHNpuz1CPxrc2avc/TnkX4ErlcT74e4bhXWAfr67g3jmU
PqsG6LK2Ex6Fxr4CtWtnBaM2k8rlH4jtlINtajc7vqe2sPginsUuh1jWiRjE4uxvJlODzOh1F7JY
naY9Gd10mSp36tSLrcNJS8+7gbxnNe0jPnD9HedKizaHUlR2DGetes9hE0Pt+nmPpUTbmMP2YkUe
NiD7CEVW+PcRSlQHU3yxqHBfBuXuWeCABNVuocoKq/LepwxhvxzBDew63hQXZGUSqAZNwfNUPcGH
4INB4TuzRONhINQlAPT7t2QlvCN/pxCSid2h8xZRGmM075Wjifc8afQ59EN28BrqqRy/qDLiPK6i
qM2Q9fRg5KL89HS5ePWaaji7nMTPZIeNJyjMQ3XRRnz8VhS0M+Hij2CGFmI80bLtqI7OpAuPqqTq
mPXPgl46C7cbUiWhU1GlyJNNq1EZ169Yb15yJ2XA/25j5uVmZN3l+0c6QVQAV/5by6IGdcWlO+Ru
OouubTuEuI+s+vRcvgiZmEuNg2QpNfZe4OBFeJOBox2GSjTkb4nNmKaeKjYkmwBOdTGxaV6R8boQ
MWyLHSQY5SZDkFpooTTQtHiF/cS1Ge7XGAz34e8DDuv55XVaxoI+sBmz23NOKQYToh51vi1sz44G
DxO1pzpo7lBKYN4yhjzsuVi534c2HouqKZqm8sZU3poloqP9jpsEpPByugQtoe4bMVMjSa1m6VPA
x8kIyQv0InrULCyJkZbdV96bzqXd40esGYACto9bs2cCkPO6HLIPyQldQCT48fBYvgJxskBj5H+V
CPxzn0xrNJREaRVzrUNbWVXSQymMouysTKOqWgYDZg8klOFpZXSe2nkAA7dnevp+c45d+XeFwOxf
Aoe01zFUCIItj2cZLbdz1OQemPnpJYBsBA6Z9ULOqWLcXe10wJp85hfcoM6VN67IEpvFSWPWKy9m
6Ip4ZYy25iPoh3Sq2ixx+kjqpFuwNRqZahkoptfZNi0ru/3eplH6gNm+ZxXdcpq4YDWpOw5ZrtkQ
lW+bCHSsg5UwfdbWs3vwiktRgquA1mPbe18lu4+XE803Kpnr6JwwTQRhgkcEk8BjiCOan8aRfrzF
cnpw70mZpcehVwXO8bMyCRzYaPUmIt8ml2uNcEOoVEXJXvG7u+Ge4ktqMjwngY64WgmAXXT7tw7t
O5iP6UoE+FXrLBT/JwEzmfD3cv91SPeZosyZkzFncNF2LoF6PpGhwdpK1SS4mPPf6bNOYmcKzENF
AzOVUSeDo8YmngxkE67cB2GcaLYdKNILAzfspQxBGovZzvVeqda/mIcksiQoQnk4RMwWlRL0LGQL
tDB853yTtEXqSVbP4XR5LMJPV2bwawvsURZNOAhExfZ6KGMcne0KX8YGIKRRm+yMTuGMxgsIIGfU
mlahnNsUVRD18G5OONUSQddPtW1rcV+DsjapPWOuHwcbBZQydMCEUr42k7ERjTvzfYeDrueaBtg9
vAbiPJDv+wMNd3xK5V9zi2vcj1ViKyjTuS9yIJY+a4wH5gsm8bMHdZocVhM9J8WFFxayse8IqaH+
8SFRBXvQ93c7c0CCCdoT77ub5x6YsRQCb9Tgn/WxIIGr7XxY727SCyMrsrnvAp22WZqUx12ODE+w
bP83cmQoC2oWxdWYZZ6SpVneoP5quEw9MkFNVRZBEyjRH0c1AObyv29o7X4e0MLfp2TW9bIT5HkE
Vq8fBZ3z5mwxPdqLf4gtjzEuWtS494bmiPjG02y5sf8K7hB6oim+Q6QImSR6f3OmoCw29+tMD53s
uvCz4rTNd7/Fq6kOmezWvt2adQDI+bQZyTQbFLvmSW/IQnOgVnj8OzBsGuoi0qsGmKm1kh/wvg3L
tuY6ZNGzygkHgOVcD4OMNLS7xfAZo1Rs5eu8S/oDrUufOWdjV2WERyyPi9msCB7keW7F6y5og0Cw
jQ6cUyJ/WPrNW2nOKoYWnAzz9HYywqHI2AtUGXcMIdiewY0VODYQ/IL29cySld6YqpfQPqKO1w8i
TDrelrILsKKCT26WQRzP2nC4DST4gy7m8zH5zTtSsVUHHQBwkv+q2DiBxrOVspSn3E7Tt9YuBhRe
C4nUtvHf8O57F02BYP39sF5TrobLObakh1dbunuSxJ9xsrjMfQH8qqC4NdAMdYXU+vY+Sm9+OpZL
CWHxSfOAupmyfzChp+9wN571IZjt/oc0RpdIjCZRs4/IeO8hvXInxJUs6L9NoPEMKPipUCF1jPpV
xV86Hf3CF8I9YSCn0r8ppMNnGwdxAHBKWLnLTdYpNF1soXHiMP+GpRuepRmEHApoPc59cW/hP8dn
m9Pqhu0t5W1QCpu1Sw8iCQLz7E8uWt+dynnPpIbdYZ5cRBhv2hbSf64WS9TRpZ6Zl5YHW5fBja9p
q9qLTzPi8chogzbnSX2owGga0InL85PPqZ2ZyTlv2PuApMhltMVM17co3PhioA8KkpykEW26+UGr
UmujiC6EiXp4W0L4NIh/XZTdsG1PrQa9sKgE5CUT+Vqu4jiUGPcS2dTW2uDrQlpbaujQFSmkElHV
5zJm/+an0m6nbVRWNUhWlPy0NaBiIMSywAlGiYZwiyAGhR9ssqXen9WChuoRVh5jEKQuG4Nj9YcZ
uZSz6vrTGhobsH73q1BX4fBaXMmDyXkWko/5RDoHNZsG+019a3Ka6mMW7mYJWCZTKxMGZdPPM+Ln
fjFBDIGJkJlUkmxFUfjwsb7xzLtRofDSkdAAyD2d0xuQAyyIsVerdAZwe1vQAOD0FZu1XhIXAY0f
a62YF6wJLA8OTMNbAKk8joHAVRX2VGGJgATB8ieuc1VCMJRu5IJ0c2Lp70xKl6poO5AI6134feZA
eqtGWASaVCty668mdFKyAy83UvkQBnp8xmI+gmcgM6UmJ7i7Q3uVauQsycLsJFFF7skl5pmqif4v
bMfjuP0meSoHg7HkfQ1pL324eVhpXbrYIo4Oxuk6taMFDEGKswJmSA3ir1Qt8LnEZH9fLZvEty+Z
Ps0suTEPog7s8+ff0zXLj6wEZw7ECIwDdbTDDvGs7EEoR2xKtOLS5+xIt4BfDyj01+jbbgj37Jq3
LcUVQpv6C/zZR6EAdz0m9wC1D1v2ZLLpyMqGCBHFfZJJwLQ89Wgd33zL3lDowSqRAP8rhbqX+YX6
qr8CCpSyAkds1fuy7e51FcutzCRRIHkhtqt9t0YYnP3Fhm0c5pT0qUirLio/0GrqdAh/hlT8MiOu
w08+17w/Kq4Jk90RP9BIc6IhE1YTG3aqtUKy+vHBmFwpaoGPlUQnV8eRMWkk2zXn6PTBmAc/tn+5
jwxYPS8nFSxpr5Rmcxj31wBHKTXjH/vGSaWo0QvnqmZ3eX4j9Ah4bJwUTI7LVp4+jKDteOYKdnw9
h5n3hxrkCiTROGdlroEiR5/ABg23WpTK1nF8aPNDStw1yf2obczj6N1l4AruUhRX4XQ5nW13fRwZ
9acz9vsO4F9tZa2YIuFPuyLl++/Ug7PdKO6/XQEZtZ7IR8oYJRoaotGJFfJwgzNxx9X2seDBlUCy
LJ/RQAtIMCg4J9QoiuZ68O1irtNVG4ZWS9Cg+ibg81IyCxW4Z+l4EGAt6TslNjArfC45XZUqqbjh
CmweeTtq3NZSJNUyVE+I+V1n2zrLxZE4V88ZeEDXYBR6zz/Q9f4usD/8ub2DyZLyvPPZD09c0TYl
QTZfm9D4eE1x4uQ7YiRDRv6qtteLaZ4CZ/fZZAnCwP1ZbdIN4WtNlTCXhklk2G5joH4ugJcG9d1P
GyIrTgIU6W5uenVNJTFbBXNXK9YTjZvlzEB+1g1jSTuKh+A2chZ18yBm92ddMu0IUGZZLc1vrcLc
qJ4u2hXuw8JldNvh6p30NNvDEnDXovpGPKKLu85R1AJwDIxZ14lPuEy0luJgb1+Etr4amfS+Iv9o
ym6EcUdZP5rq1D5BYLBRUgn+nU6GcgkiHtZ3PXpJj4O1m4YZOBncLBucYuGnQ7OLrLh88aV4lx0H
mzTrfSRyUism3pFH3OWOcf88/TPf9iSH+1QqGqSns+vDKtUss0vPZ06KtYVw2GHRN+goOUS6vtOT
IKmEZ2SmoZX46+CDdaehTZPVqLQBvKt8+mMPxdAUa0eYICJ3k0ICa1uMmWBBQN/36rxIZyH8EmIv
r6tWeAfOEZnhuk3DYmKI6J3+xn5jNHFI3MCArZTTMb5qBMtftPoYxO6mJ5Z1GVZUPx4K7yu6lKLZ
wz0uUpP8ecDn9aMsnPG65mYdWmeOviRC1miCsXhou5csvnXEvTqJnMiWEuEL+Sjv75Sg+wpXyRsU
BzU1kohuGjwDhOXL+pVjl6NxOvq1RYVXfNdut3ikkP5x+IRLlhSHfxqBr+cRVz+Rbsw4u7J8XJmI
9qv1CKuEE6f9kE+15C7j94Ndop/7T5uCNec4i7lvKyuGxRf3YAaWcIrD6t0/kw7eUuHlqosFwjoC
sci9xcbpJGQIblZ3++ZB+iSq7pAAk+1+XehMFD5zKJGMl6VE7JiHmwFl1HDbIWcspN2qDtj5KfST
DrJ3Ev4DprYx7swWsj9VDqiwmz8q/Tkj07g4ytQofUULoTDwhZ+TFgEVQO7b0hViTcuxfq2fs8Hl
zBYq2oXcBxmHTj/Ef5qVPR+SjtOTAhswQxHc4ixIyHK7xQWzf9tbb4fje3bDqREV+86lQOfdpdSF
VKHU76ykkH0FOROPGfeSyclT0OpVoyHnCoKxJjfV4ShiVLrS8etKmLFIW2rLgj7VPXGHrPLQwMmI
55fy3l+wWmgzs1EiVkxytSd5AqlHXgEwNJYuMoQIa51iZ/LIvKTsYf4Mw8JtRy6vXGpmlE/65ohN
yiy4L+e5qETDSPLEM8+NrOSZS91jzCW6K0jMaKoFJGrnTl2SV3s4W9yxzJ9nVx68qH19JxwP8Zfe
+3bhtcL3fqsR7lutyLjNJeKZYIwOJVx11Lr78L3swMucBL5W+WNrwg79u1wp/7qr6MRThuWWRike
p7myEjf3QDoVqr7+zr3A4DhMbN1CovMDYsagpHXxQ+qQyKSYq4m2ax8FmlT7Nd35FC4n3KXFz9br
7ksNC6ozpP/T7/MNRMoam6HxT5eeP16WfVavuAZ/a4JiZyHGyixBE0XRkNINt9UIAAoItEBykrBf
CJes/7dd4oFcyT8UpFFAYaPOfQ1F9UtBX/Dg4AGO2Yh5kw3muUJIc1mv378kYy9+CgtXHDOcV3D9
yjwrtVXZEefClFA5MWWOFrhyL1hsZY4XbHyVo7Mc/+NHL0D8jj6M4WbcsjOvl6hw57Xm8KIN0gPJ
EnE82eaA0n2DnIhaRzI/C4qKS1IxgWqwwMuGRIzKoNFV7brrratlhX/TbyijzS/3JWoK3Bm1TfUk
CKtxWwCwGdRUle7Egi3cYFD14ArN9yUBL0zw0ky+cSKub/Wl/Vlxy1u6ouiK3hmvXF5ttNXHXGm2
wnqQn1O0lfegc3lRaSo6OMDzjyIs3St5KSuFRk8+j2RBCNOtfNlyGTihhh3mWk5Ep+7uDnJnWw7m
6dq6IXlPWx8zYkYd1AGHwAIXsiMCYnR5QVv4L0ShhQF7MQQshxX/VDO2LecdAuMcs2l5njQwuL8E
nydMTKUMJ9f+08KYJLsJZBSNfblAE9FdxmcsOFNoQ8PnnJdiKgq5cyNgqtpbGHmU4mt0Fn+gCKLm
In/3MkMcxpt4qRAhKpZXH+AZJByaIxN044DOf7enR0FQGkIveN6Q4ThBQb8LsEWJjDOVtLN/gu0U
eMHDObrt8+bSDH8e69hn+SjXVXu00cauaCSs97+PeMhFYBARcgWruuj4Zr1MqlKJLkDSDrz9LIF5
W3nMRDgvFjDZk6I8845fxNsTyztNyNXJpoz1g3icaYatdQ0v2siaYBwBfzDEDT/nVdW5ym7NlYk8
zOZSE2vjGLQloySWwjFDmNYwGp7LdfC2yMxmvREsxCSTwodeUDH02gFWCrfOXuE3ShyEqJDauip1
a9GhKmXuB4ln3LgOWMYIFJkkEu3G//ERSwp8OHiS2/xf/JBnoDjxIDCmJrQA3R9lCuhDMxI2feQE
zfEjMREap65dS8xXGqmsuMIPV0V9bmhkdCefVCpdT1JG3BZ45WgPYm1e49tNZWfnbZu1AHlXh4HF
gRzOsmQ5mt9LgKUscDfvkMYuD5N2hANuetRBV6gjygREWxt7eZI0GxFtyvguuQlMugOmSayHljzw
WKieIKydYb0qnieiEMbyGxZOIJDpAmA+lA5hDBj0Oem0sIulNEBbO0EvkLCSZXgG0X3j6UhPBm3O
daEnPVodc9r63OjyqfUuyHFDa3EENjKoT4xPoFf1lElCJmo8RpCf4i9IZxF9NvI07wc7oCoGgrEy
nJuGqtBzBiqx9K+H55x043iUJG8yLO0fjikiE73xiX5G77QWUkr7pUBNndIkzir3otr/cLlPdeMz
rjqtisS1T944JpV0qwinKhDmZvQlIFb+9u2ktol/i3CVh28Yj8m7zPsdMWtdavuqeZyUuaE6XzH9
GIR4FxQBhO7HXNypqsG8Fp/1Z92NCijSSo9YkWdeGe5xPIKSBlFJYH2UtR4+9plQCLLByVpu5mGy
Ag0RVwMXmFW9G4G+Y/YK+I2zTKymJszTsRvGnIDFHHM5teApqYovmC2v1IzjZyi8Dg6Mz3Tzvki4
aLrzsQUC94+1ERbD6crOWKdwsXMta0N9AX6ZDnHhc73G6t5xgnTZv97F1Qmdpw48CmfssPseFo0Y
B5IoF2TFmQ/AE3+V2lQN6S0oNIbqnVqu9en7cpvZG5D6oWwncN5tW+3lopvKmwyYuiGRnq61a+bo
Yo/4hTW0DXuROomsj6TMoKUeshUL+wfVbirDzOnZRjI6dDo6yk/ZbUpSjva73RDzyqgcVegtBFDq
h/HCqlDoPGcOMVTdN0IWujJw+BEcFHhPvjn5WfLyj8STpRmCeAFT+PA11JZ2OJgFOwgEqiuXkBZv
3ZELovElOox77tqI3vlfEgWUut1GVwW6KT89mYd8FvZ76PzgO6EaNboUxFXZSh4Sc/ccFIN6wf+v
drMKXh+TfNIb6J9clEhhIAtyCsbmO2NMHKWyZI4ngc/yOb/OeHwi0vdIusBkB29TYzsQ1oF7VNYv
MTo1VYta+PtlE03ZGftGD4T4uWasEPGrGIPpJYkVmOCBSA/5pmPhsB4npQVWdMl+gH3XniM2MpUC
L2ltnOWFiu6bPfhj7JXnQk+XdGovQ1GnCd0rqo9gjSMI0y5y/LSnj+wdTsorUD03MAQZdhPeAGk+
CwBKJiALkNdAWMh6X2+G97CLnNgXTnGMwNeas1yq0Bt8RUt/7Ktwi+BNsiU70ZSpb5urGxjL/2Sr
CY0g7tCWkFVgM69eOCbYed8bZyKOvO32DgoPZ2JW4TPnGiQKDuma5zZgu2fXkAEPpNSFN6fN0cAC
AJUSM8ngbppaRHDyqzeRLir8MAIx2yAaTTsgT+gL7bXvfHo2dIyMrHBcoiupPnhfafgKjKeMdC7I
yMfk4MFHcrc88TVfEV9UlGRkpIo0qFTRFMP59YV5klQGiogjfjOc7MRZf4BzoinA73uaYjHesEmW
mRdIUP0/7cWgoGT4dF3UFiqgOUC6xmeCG/fEVCDHWvsyn9Bu74fURbYGO6R0tRP2WN0lNiVHzyDK
fCqwnyne9pOTPfbtDsSFJnZp2TtPAiJ8qgqojRGAFQdzCi2pEJSRrlJoALKDY2NSRLVuVSdcutRf
ucOyu8W+AkucW40nYRi23x95wMQVM4/9DE2YNyZdCL4M+xAzDBmukJiLGXK6ifxrGKpplJuwR9OL
5L8pPwi5SxdWKvVGX5YtCATweMNXlxa7wWx9b9EHKcUWHg6E1OzWk4JW1YRji+5ZoX31RinOy9SQ
yMPz6KOlnlEcVghWjOKcvO6bCyO59BcXWx3JWFcbIHUmOfYsOL9VPJcOuSYhDpSn3Mau/kfOwoB3
Oscd2YMeRHl7LK+72s6gxTYwirBaqHOnjtHN/Bnz/EOnblfkLL9Cu35N1FL25gI+yxb0VpE05SfA
IeapZZ8yAhIp2c6F8lHkLYaChCgKHEqQgaigoBPhzRa9LnjFzXvSfNkVvw833kiYEAktk1XLzhcP
zklwl3sTjF2ZM1/dAPxpXEKlF4n5/KOzIoUsdRGteNMiwhjYr+F6y/l8eKMHSc1LwUxdOkVOso4o
Fw2dxCfUg0Kydl1w2MPIjNUdftC/GdPoIw3YrgpiWldPQUDgcqIC+lRqbyiIr5ETQNSvgF9mx+AE
l8yW2ZprqlGfS202bl7Vl8OMtxynVDg5txbTqUaphuSNCy6j6wUudyokRyfyyRgoO5APyUG10SY9
6MWSrxxvcpG444OMv6YlRJxfHgjjghpMQolK5adTOzC3QRpF8N0mtb2TV5qK6jx1Tre0Rfqf26X3
SmWv1IE4SnH5a1t6fsXVSSu+gVxvGYbBpH5rR/nVtQGGQ8z0NNgp+C0y/4C1PCBYI6zCYCX9alTI
07lWXhMnXkzcEb0pomuyRoOZXZPMBXRsIbQgi5XdWLgBSjaaHmB1NxJW0zj+eRcS/5Nyktacr7Go
PtPhEbHTnibD4Qe7YnC9bYCrupJyHU+ZmZsOnqmsd+UfUcMJxYvc5DpsGVBrpIeYIjew3C84+ZiA
pGqkedGFV6LOflfQpJgMF0EymCUdPkAi81deYo79YqPp87PMtEPBAKGGZSWXluOVsyh2WB6NRtd/
ewl5cJOAod36cdlZ1Y3EXyu4ST7QnIvvOJTbuyzfvTV6ILpMSNplcgq7zncNxL/dLAt0G8nRRhwt
Ov/Rkr3YddXoxlVfNvNrEfinxfvkFVmAp/TLpS2yew4KSouoHXUjyvEWTpmVLyitmQOoXrRFkg6T
lpXqXPrMMKJ+tU53ERV9qK6XCo9Y8VV1S8K1AHxDRQX+DyiJW5mJqLga3jbMbGTtKMOObk+PYWFB
oBdIgFgeUslLzonXtyZosRM7gO9MjnWyXwxDI6UG/U6BZaxB+4tmJUzZNthwyEt86b6HtDE3IuFW
EP7pjCo4fH/kc2+8wNM7QquM9MlZTjQC8FdztUCHg6gjoYQYg2Pa+cXMl3UN4f97faPALs68jPA+
Go8ymkNaWInEkYSSBT7GvZNVX7RLDLvrrGpMx8S+iHYjocjvF4WhlGYYFdqkGPuBMnF23fnzqgo4
mw0PQ02LV5GTLwWVuSCujMNYyDXN8l91jRuHL4belDcZPh1Ss8CMvkArVX17RUzd1EupwHwXweZk
YzYYVtOLqUodiHyVbRvz80nelO+r1PfqNGtyFUZ4vxsZz4LZ9gWKAJDUEkNI7mXHk8FiZmSVvHf4
B/Oxj68mXRyEE4zDbLvLjkRv+nlL+CLigZV5uDVO/iPeE+XfSoaXAVhSBAuCSX5ysHJ7nmrQeF+g
BR9sak5p/FShU6UgK2xeIfKHTWI+vCQbbTINCApqyt5j0gHcL6cVpN1Jj37EVJDfWhlb8PI00mRK
/MwpoB5XctL8ctlCSaJHHD36Acihx1fX2F0VFYEoOO/I5lVESThEvaEBhUxBAsK1aVAWPyqYjC1L
qXoiHVfXVG67kLp9/O7Sm/mRvbL69Lnkvq3CtbeOLkzUpwGYT6eBTNWu3PzfH/kTRiZVS1YcKTSw
hwfYXMEmjcwYx0Y35tFZZehNdx+OSljGA1E7hDmrFxiHiPmYoeCl0T+bdMFmtRkZsDSyErJEpORJ
JVQYjgGBnmAqJUKjhBDTAfr4BbECj4o6DSNPmo/bSpv7KAc73flyOJf4Ijk+hQ36m/mAq7H/mu80
Io8vW0N5TqrzV3tmtBqf1njV9NXxKL9ZuLNDc91JkibZ4Hj+31dAWalcONdB0zbGNGbgfZaWQgTV
J+eLJlZhgcj8Y8R06fJwAGNsvTdEs5IwQVQfDHrJzYwwlLsDw4kfSMo7UxU7ur8EWaxmfr9VOWM9
M+9hg0VAjkhm1QdaUS+lK8/hFghFzvSqeI9dwo38DOuEuDLUasVQ3LCMVMfACggUDUSTC0igEn05
uwzoKZLIWC2cMkmrhu2poQ9NOwe6OftCHmiW2OxEHOIRd0AiBDwz8Ig1XrxwvEWVlIhzhWJC0F66
c9/W9DpO/khA/fiWbgds9bMXcJxo4SaciB/UrAQbhr11+NHfm7Y3KikQWojN0esKUUIB4GgHSIaK
OYauhtGSk3n1wgPuARQbUStqMOSpHKyTvv2qfelu1PsdNNvpLKL0v5B1OjZjyPsyv+vhe0QPfaNM
V+ppi87V4s/+ERH8cosFKdne+o4rLjmVUbFbB8sRz92UE1ofd90WSiQ4Gu4OdLQIUokrQ/0WYBiU
HkMlL7/+oEjzk7Ur/3sUD3BkGJfuxZxX1XQsqjFkVCyc3DZ8rXy8eMYHgkETBXT8QGLzLnFLqe3i
kTBiijSPjhbQZp3zs1GByDL0zg/LsxQjuM/FTKH7c8zvZvOza1uGvtb8l3mq53+NLCGhIhr6slEM
bWmmLwR8tFKNufq/KJtmVRAcUaMw0AUStYYb92Iyfdxkj6EHM6v3tclrZiHg4AGDk3Y2SS4yT7cA
jHRnhbwMCngTV/PaGwFdWCQRFCLP1X430Gfs0XFPOykTXNCWTYJG5jMcyQ7t1eRobimb2jmNCMYx
oK0cHPWf0u8Paw9vqR4So3p3r5bSoyH0kkwgfjf2ex2wrmh7kAiCD2EIk0t2BtRj2JYt3aiybrh3
1g9HVBcOpvNjygBTblHIsLDPSTKWTzBUEvpORVZy14WEYfmVc96mZrgoqFfZUtbDAgf0vWSXL+zB
0GlkdL1urEMdB2hsacHT8elEzXjdpgSpkaIba3lIInfUbNxYJT+/erRxN+ObeVZSGVr9kb5AUsQ3
nWomijBwHQkd1S2ThMmahBIA4bfGcNgRzjMbtcmyJxJz7MWZHG7e+ABHocHVFqGpxgRys1Xlwjlb
/e5Rw5gFnc8Caw2lECHbIYb9xcbpuvyCIPKMMUEHZIXb2zTF3xYb1tmvx7EjnrkhOeKbUNilOjkF
QoemR5B+5dRW+XXIiBkxK35YRLeNNbc0Pe5TKEvP58mCVmdrfjYcoWadFVMKGCiG/1OqqIHd0W2a
DSDDFkz1GejuFIIzcH08zRwdZ4K7xwv6Gv+OwKf1vk2favyxbtqOONimcoOGLfYQzf/sToIb4D3x
DpXGmJgJa379MyK1bIEAKqn12K4Qtch7d9wMrxh+O4U+5e1SHaLn5zgdts6bhH2Up8oEpw72X7qQ
0qe8hy82inecndiscCy1zGit2aypLWshUNFTun0pspgEzBf3kS5EkEXJO+SZBRqgq0gQCCPp2AV9
0SWdSM7GQMdifeqkR0hRpkfX8v3CWCh4MBIOzuBzgCOHukzKaccTUbnu7FiGFvIKuEneRRuD6m1d
o3qdaqpubFRcZcfH8QUWorfmfKHZVGDwxfEpG2i66763/r8fQKw3Rgrcw75WC3p64rDF3tr3P96G
n++Ga83Ql1/Qx1UPwdvMGLrho2UtbFJL5lifCy3b2egG7wbkT9OUpmuqNOPBylzSZkjrB25E7M4y
qnt35UK+XJuEghYOPWwv5UaZJi3tTE+JOU6m26tL0ebigjPfgq8Z7kHUkw9uomdhfvVlXmNOS4fK
eodYhIqZzelon9ZTcFCZ7PA6g8wBw1ilysY3LK8S82M56loQ9mIw3SxFy4erD47irpxdco3W1ZvX
QFa5ulUrmCRWsy3V/olefLeVzt/B2qZqrk0lgFAGWWVAnbw69IsKjkweEETV1TGJU1885p7ngLDe
tXf2r6P4po8/GMnctCq8LHRtkoBAvQapoSeyCsEjuAuiLHDnGQaEzN6j4y0Mp8jLm3PCW2IYW/8I
P8LF4zxGQGjdyqXvpFHMB1B7LoJS/lh1UgLNnbiBrJK99zbom0XlCpaxER/JcfuLkb4SwLF4ykmy
CTTKze8n2j0XdUeIhy3ffluJCY8T4lNLZNEZJM0qGpBVAaQXCQ/cuwdrHwhcHCsKl+hIbmoHTTnO
SuqFKxQ6M8wBanLW/oosU0RrmgzUvHtLINKYP9bbk3+Naz2leJ8+ixQTVPltiyPyDUn4+S0i0DZB
qrPdZ3WnbKBaDn/YvteyGRBDuVfqxBnuMJlqIQGnNaVpLJVEBV8r11zgispL44Y9uxWXlI10D/iT
Fbr8g70eVOn4y+6nvkLg+Ax+i7raSOCFXsXm934LIECfKpPXeZCCM474DSSTUlJDg9aWwPcT3VMM
7vBm8D03GBX0UjaVcffVpcNRbw3p5ZoQXgd9sSVa4l/FIfRAFbDz+7+FBmy04ahFFVGuJEh74b2p
6typkqUIxOUL+MdYOcQt5ts00yx5Z8rl017gaMUedqCnB45XFV4eYVsnME/OsUccZbk4dHdxa9i7
wpftM7wrdXfx8tZ7fYpVZYgIL34iF+Dv5wyli/s0+znl2jyFfhdncHhyao4zxEGYq7Ai7+GZTpiX
pM7a6k+wTFQVjYUAQ1tTjVTj4+rdAUDTPwS+72rwi3Fe0XSiswrT4Xui8asipEWq065/Z/YFFu67
gXgJyyTjNgxBhBDxySmeB7eP1LjuGAbyir/LR4cssAyxWP/MosXu2rHpohcdrsONVjzCq2+41kx+
O7PYwh7OSIP1y6ypTtZQtK43+fM/0s09uG/fxNqmsTZHW1AgqjM/N+TuoZ7Oo2pwko43OtGIt7Pr
mZ0UAR1W3++iz9K8Fa3Hq/bRcGlhbB8PHH+hTv0J/Pkvjk/TRhMONh/5qWP7089ah1mvdMjAz2mo
9jmCNBAwVhIgPfVxGkJNm+R8csg2WbZ1R9Yw3GG541uD+pnVKs5VhY5ssLH11KD77j82L1UEh6RT
fuPlZmxd8BAXlp2wZQhyDJom926znm+3ctasonwxxcYioX73D8LqkZdix1vaK/H9FSY3n8NjncbO
fPqoYChPqhZ7LNIQWHstGlH1aRjpMxOYDgQ/Mc1oplTz5mlrqYU1c1O091jG723OIPSiEQikuBJG
d2CikqfLgcIZOthGtW9J0kjKBEwAk+nrBJXjZgaUYYprAeSwYiGi4/QoJmN0bFFm/Qel2dPvI/ZK
oiUee/7a2kpJz4PbUpJdqtj/EwYlRYU5f1UzjpXz7n1VYKJnUTm+dv339WZt1484ksAH2pwIIauQ
VfvbXyt+hUzPha4srl1BFiIF1LroJ08enxdXkkqm2p7fuMWNBYZXVX3lmiGpd115E1FEhnZQ3x57
EkW1DSQwPY/qoUMeNhtPOjEn/1WivISU+WctMsoE/J1mNI4tqV3Hmi/nfmaQI+T3bZOzpgbzjvrR
B335eUgm3Jo7+db/Re+l1hc3e32wA/anqzUgwj3SRc2FWcrAo++YW8c9FA/200wZ/JgBNXuAbFhz
lcxkERLJWyvUNgh0ncSC6ZoKCFbdriecmbiKfPYgXznS2Iv0geUoyWdY9DUHmYMHL3frN+jL02oh
2N9PNY5Vcq5s4ebJFGsOJWeS0WTVpkASnC8WvreOoOFr6p5eLCNMjpL09D0HcUJHWx/iYlfp30MS
vuqNa0IVO1+b2sDoLOZQXjVdL/FIXmWWtZiJIrK9zpmNa6VMW9+PSgHyp4vaDiHYsN8wQfHZPLrx
jO3ngftrjnfNRbXuJo4sfCUxZeiDW3Nw09bCPhTcntSN1B3YsB88lZ4aacSI6zdi/YAauz6sKkCw
oGpgwGzZM1NUa3mVijwjK6rx0Z8GF38tNuji5i02vdVVjvedhA2qTyMmLKpzsuuZbCOQ5+dQmqv5
1WfLPdIhfbjWUZRzb0lYPG2/+s2wL3kBa/pazSR1VENo2YqW1obmUPHKYeHbOzAnUIZHjEA8N6wN
pkaMb3d5Xi51EXsK8QynoNn7iWEkywTlM5Wa6msBMf2fsfolQPhtjnSb8Vlfsa2856M0M87oNttb
sXnwQ0zYjsjpgmI8IWvVJPLRFhS8DoY3j9byM0G1iLxKrTXuqtDe5p/QTzrvykwgOEQ1ae2tR5RU
gzSwzqTb/MFCggUvKokTMXAZDRzr0mPEKJvQ4skb9ActFXGKGlaPlOmIXy0alyaVDcTEQ77EcwBf
il/Z2NM5sUti8p1zO1gU4wtPq42Ocy28R6iVrmxqH0DP/1sXivpv8D7zEQV+I0NtbPcLE4rpGtog
tHtEl3YhRu/jvh4D8pfPNJ0I/IF+QePqXcwLzd9xARisx4jngrB4cBpse137WUEluXnGSsArjlZ0
xCzQuYLcGWgrbpEXcs4FdiurgDNhQrHY+n1yNWa5y26bB5Iq2F6sVj+1zt5jCQNs+Na9qG8PtDl8
ak9JX/XLVrcqV0Rt1RKT2Uoph3Onl820UVOpi3VoPtahVuCX2X+T78j+sXb+IECjR/CymhV88jBe
Leg9116JO9LM4kW1+2RB3NW143FrRyvbA4Q2ImpAdSJJ0niUbMxmamkGVgEOlhAKw+rv4Gn2+yPX
8/maDbDRbnQXVpwbiNBKLvPyynW9W7sdfN3BWVxSmKb07oz85eQs3UvcuWK4uqwrmFFs5dEBFoYZ
vWWbPiHBQaUavd9f20uOPlXEaFnU9dNuEnvYHEt4Mzy3agysqxUzsv/UzGy4r+Qmmz/LFS8NrNSn
+/jrQ/kc/fzYUzNV9Z95+h3l1d+Id9BMMoIQI303AoPT27ovg6wPlp0kE/Y7QiBI4/k0FTOzYP6W
5iglpqmh2G2kmJjdqpol569NErz3WljXmactyBw8mv1aSzs3jWz1LSrvx706nuY3K3FafUjb9I3y
7taRYhbK62xawM9Ty2wipFzOCbdVLgM2Hu3nE3FPuCyMVDxMuhUVIKr+eELlX0o+/JirWJtBZXiZ
fhWaJApnq4A0WS5HgTjOZUO66DaMAUsiNgNyb+YhGPu67lib1Jceee56ru/1A2+A4W78Cz5wxjMU
fHJfdbazrz/U6M+2CauIHG6I49UU+qGOrBDgi8eg6nZMuweg6ifyc/6GmESn1loH1RQtz2MtGB3D
FEvmrJ2rQqx3KAXHVdIZl54OoJsCSQ2Dk2D8OKD6YYApNR4oBQxgEmmCQOyCqidz39ldqc/S+DcX
h5/iJRjQJj4Bs6XY8rwKZScD6q95juNs6c1qJyt4bsSGMvQMC/MqUI1EjLvJz6fG5vPWeAB4jHcO
yygp+URrCtV1Mi7PVccBMTRtl+MsmqiYBPtmN2OXgW4JniUMg9ZEU11SPndHRhjeyAlXgV9uGpGw
Gqft5g6OujD/7pc2iew1Pq7aG8ie7zSiuwhxh2USE0xJ0fFkgrZTnPDKP/8BNG/zTMg5AcSb5J/I
UY+Jksb0LQwNQP+deBm+dXo2fQ9uYdvO7LYfuVNZ4+vDhX5TlcELykS+lOUg9ajTYwuOoSgYC0MX
Ld70BJNkByv38f9xN0KhFpEvFrw5j3vgwaSoocddkw1jAUEBXHNsM+WEnUMZbXnzYzVcXi7z/ede
BIx2ROvr4suhaeNSBxcjOSLGXp9MFHzxnyZwETzNGVtRSgQL0UXc7kueQqypE3SeMucTKYTu7AzC
XFkIXus4TtuqIDq8XI2RsjbXGk1cKf6k0A7oDqbPMs2E6Jti/Sq+iTV8A+IDQS80GiqPyrOjvFnr
PT7si0Pwq6HPki4sVonkkyuLqqYLgwsmE1IHO6cPcTl9zK6htWcu74XD2l4NJoJA8kMAR1XI/6MR
JS92gcul2tFuXuY0w7G9IRIeYoO0NelEVpArdrawkwi7pj+biev2h9Ky2z340nsGqNhvm9DSQj58
WTqoSCMlxNvKLDCLc0y1t8Pb52/3aDdKBW/zVyZaP2YIa/vfDayektdhKkuGGc+CWK1Jqes/A8Jg
ZdIT4nmn6UjAHPRWpnT0ZrWo/vd43qWpUK1jHxwTwNqkljQ6hG69psPZA9mQfUyuTE/wD8zLQ0HW
I4o7ZgrUIcY/6H7N4QWHnOI2FA4eoxH4NpLomQ20rppt5gFRPzZIz2dTEpMi69GeBlB2k4Km8plf
0EVezbgUg9W0SOzbvsIcSUF/Cfp+9jIGFodEFGDtzp9Mxlpf9vO8A3PqEvQ2o+rOSc9J49HmPubP
4OnBxu63pN9b26LJRyQ1G+SsV9tLBYEBGKrsh5SSF1zYL6NwdAMqLjhiZ+1OlYWAw5fdrnaN75tb
c09nJ69HqhZkO7cn3KEgEiMEp6i2Kl0ohddyL7UV0FnOHh3EEpsdY4lG3TrrA6StEr7Q3hP6Q+CX
EggP/B9IsgZVAx5xZ13N+KyQsN3ZBZm8txGtIF2x6Ch0bgeobQafXBvMJghufZEd2SdOQY1N6raF
y13gaK/sdK8ksD/opJm1v6UAV+pynCAWB3UqpP+6M7GBA/8FBJ2AEL++PjKGHm0RSQ5lQ686ah2K
LKeSTgw0r1hqZgwtj2dkOk/LHOpeRHDC841BABpCnwRVvRWuVLJeUrVn1V6JjrpAglgwDlq6XvM0
w8my0qUUh7ryoznir+y/xIw7tT/FLvot7SS+H2l0kcQIob9GU2wINo2aFgRJB9yWKp+Fcepv1I37
7VQGArdM09b3fWhNiB0nU0xrlG9gddjQk3QiPF4+BUWfcDRxzF4rXt5US8MyCLc0sPMhbJcmguHi
vCYHzh3/TWiH50rHvfpbYK64qa1Le4+buhcw4nGB/xqrSPeURgvuovaYrJtMBo4gyo51vQBq2QBp
JGwiETVFaC5HWgLpAYwbsfIuYqsqKLOkI2gk22Sj07tFuznffqZS5JWhxLIqL9gKpiJufYXxpa1g
Hoa+CgNJ8/zk1jjJw3JV/cBv2+b3oSuJyXbRGnpZ37NA/Yh2cK13nUEILAJmO2yT2Z8QGoJnrADw
ff/c5uLlxZu4zsPgU3zmTmmBygfaXeL47cdo31yPT1Rt0UH7pzAcbs+ITBj1s3ITqcM2GIOgt9EV
x7SUjD4QmcOiPjjbE4yAr3IA7gib/s3YKBKpBoJurpkIYai6jl0vdmPhvtNAFvtQImxMxGRg8fzv
mWj95vfJzf3KNLcWun6W0mVD+7G9RfBDY/nUoBIZe2WXIat2gck/JGBAdNgjTIXWA3vyM50X27yi
52hYFBLEY9SzoV3uumb1fLHN9AC4GNlWBwfNaEAWlAYEK1AfIamMbl7dCrjGnM79ubVBDnAQzULz
o8C7Wx3XH8Y0xMeklb81ZJ7ivX2JBsQAfGvfM/UzoUMZKTRfQGwPCkH7dTi/owP+hcPDp65BAvda
YAJWvs95UF/JxjFbAnpxQa2QEW2e55Gm3zzzKDSgNup3U7r3TtRFQx9iA/0XYNOmqMAzbpumBLD2
IxJax7jCaQbfh2S/mdvFIyIJR48nfpmPDeHEJOjNuhSRg+EzO+IhuylzS9bjPLtioEyUNG4J0aRb
umzt2LgLmXRwp6l1MWey6FzjclzAdtI4ShqLefCUrWhia89dTwJZqNcrOHzQcBStPtKXe57Do0ci
yU/Km5JemlmwmtfmUeal4xC/STLuzFwe8lJfYP6HXAokvZmVtxIuHN23aQgTf0atDOywONYmPSqr
7IZth8Y9WTGt+f4yT2fNYu/Z4aslOFIpO+TSUUUVNrSwBMXugyWDn0tpJi4dtPk2KtWCOYNgeTgw
Z4j5GI+kKv1GHyzohQ4BOzwbX957DWsiZgSQxxzQEKs0KKLvYcUD2gnZm+lPG+yWnbM0nAkfia3g
Zt1JKjWEwR1ExnOi86m9wsC5nW6K98K+CrGGBeXCFyyNQOqUEq1SRZDHPqh+hci81HpHKlaTnWBD
oEq6tz+ex2U85TBV93GBzyO0jbFiQEjpv0liSfmQNYbBJL4OMIbbub8k7I4WmovthJKZ4rlaFY/8
xImcih4W8ud4v/5BeIzCMLNqsBrkExh4Zt8fN1xew2pszcohKHgOsh3VJ9TmVM2ahKiQruJaUH93
KR/+sGT6vytfVulrx0eB+X2bx2TJls1hbIMp267iVLNHX6S7uZOCHAK2nFjZ/C5o2yeHbnGoNDvi
vvaSm0eg8XAcik+O9k07BuFoBIuaGrIOBedJzX8DjP9kb7BcLRuSNaWBM0Sx936IXWfT9rwJcxmZ
+V9faOC/zN2CwaKFAu3YEoE+xvA3zZ/ubfUCTBKNtcvpfXSN+QLZnkjUPEj19a0padFSqpyf6k+T
gKgy4CFinlDMc9Xv+6eZIODvzPe98pwXmbKiqlRvDca9g44XA+JWZIh5OMXNRlP7nYq2nW/VW4Ax
wX+yMcBOUuS2L7nXamKcx1aO24rHQeAmfj5wxF8duAqjHXsW+l86gEwpM4EXZ2S22uiib+cAlLgi
WEZeDEZGWA17MlLV9YpbDTpjRnmiVgIDAwRJn0988FVNGUbt9lO9b/ncoUXSqK59s8ZfPKZ81Enf
lTmKwjMlTDJmVhH8sdw/kEC9d3PtJ8Aks5I4lsYcBQVhOQq3zxqNX8EvIt5/T4+xy3c160DZqImP
bsLLCk2NN2YRCBs5Dp1itZa0MJfuuMGvFyHQ1w29/HJmDj0wlP0BnBDAzm3AIG3wJOFY64Dp0Xq2
WbhuT25gVq7yQR5eSApUQcKp/1SKplskM+xO2GAoj9qJup6OcLcgwhK5p8A0L4f7IQaQarP7awK1
KrJ78kGRIZ4x2aDp3RPpZ8AZJqrHVWvdWR66vqpbmveuKrdbhTogBdkrwxoy/DVhEPxPDINOftq8
Lf9KTfc8dudD/K3v3OSMefdwN2KbcNHEut3biLmdwhoDMCtbAkVbbAkwOy/NxMyxd0kQMYU6r8Gb
NqgpQRmnipFPNRU/hvJMYLuqiQv9JNEunkipWxNwDUs1kIBkxgEiqx775td9CUL2WnE42H8K4uJE
HX+2QPahVYEDBVgoyi692TdYOEWh8sIhR2t+EaVn3fGBV1jyMNGlcf6SaLtKMdLROWIFzmqAXV5z
896ftx27Q1V4MnoxZPiDY1loLXV3H9fvMqACZSz8T1BYPTlLOC/35RlRyQ4nKHwuPAJ6t0/KcEvX
XjlhVM278PT8khxjgdybhsRxrE4F2SfnAfDC0wV60+poFOPtseuEZPfVi080u1HSlEjR2LfaF6ya
U4I1QkyrpOge/5ifugPrtTiagwrXF0yBkmOpd3B7T0QonJBuJv8TFbNpSAjkY5jVdchdo1vk7jWV
ydJb6STUJQvM4vxCH2T7eBzXtrIzn9lnpsqMDi2s8SmH0myD6euWVsMSpsLbPNcNlkFdLAQSsrNf
87Hx9Er4nP/qsKyktr+LyXxke8VUpDrP33zGorDyTeaCc1ejQBXLqmI5AX6IGoBhGXV4+fR6sPxe
BJ9G/SxfY6N//2l/nzbR7Hc98ZOW2VYy0fknRP2JeB55pAdgxgCUEaobriT/dXN2YF0eTMHAqhXd
qM9KG21gbKy4EIZ1we4KTZnzf1d8qe0tGvx7Ca4T92aYrWMssEwnQSpCkuygtNjNRJix2sI4IsV9
UtYsbiF1ou1MNF1A+sVkQFj5LD7oBcoHVPuDUvzmA/GCVh5ZCcdok0w12atp1xOgiMbRgEKPykak
7VGFKjEMM1XF6M3Yq6+7g2umFSPHcJCa9NL1a7LoGSj650JuR3Us9k8+PQzfDIikcdP1vUtVsurR
+msrb814iZymJk1N5i66i8WN9QCAG2tSxRuAZed2PjCxQeoZEUH4OWEi5jUNvOnAzr9qjea7/no6
Vvp2MAPoOzSvEh2T4IpHu2dcBNU6Q9VGAEKRA0bACYFSheBlz790bbb8ikfFS41mqYq8xC1bagD+
DjCMQ11xAeBPT43MW+uwEqsMLl0qRt/Q4c5jNojr36TINvZy6jWv8GzE0qsvqTEMHTgZY1DWQ0CW
QN+lCqoGxdcPShnsPrqQsQ1Ok40groRoQ8Aoq53XEerAXCXV6/21nTiiS7s4OEPDi13yfbj+y/5A
EmfDGF20Hti8D9DyHC+ydi/Q6L82c9PgCfpCDTcENUh7xiijUWgeoykZGGX28h8bVR/0hW9eog6q
5dEKmyPyxw8a5X8KoynFe/FAFA/WkYgXT6kLhJ032Ej7HsDBz3ANJD2GFpDB1etTPGpL0Vj9qfiO
NMlvkeTZ+C1q6N8vhmxKKx1y6/nfiAI7BPJsU2Ceor1f2O3Oz/7Nr5NZiAnWy+py+Bd2Grpw1Roh
/8z1nEGF2pEZd8uElr7euvx+rVx0QePA5yNDyuTDvt4wHOhEQi48JVI7YXAoVgtjW0R/JKkg5iMm
J5fD6uMXqc2WSCx3N72Dk1gtxFyudsRbqJ/N5AoSKuaCYg2MxKD68AzzsTb9zWG5oMOGnFyf90eD
3prg/PVZUc7nmnhYso3X6T2r27qq0ssKMd/+UootM0cl7wDGItdbz8/vh65iyO0WAUNWpdECQR3E
wM+VgqK1isKonTG85SqOQXWoH+R8p1CCYHfGBhS34RYV6YHHlafxehzNRHfvkLkhbbVAUmOTWR6r
NR2Ch21Pq7tuH9yiUu4HkioDMhv63ITRL725yn1SOpio5GtnqVNvSz76bkxXjHTVZburu2wgpFFV
asHUoPltc+SYKmig7Qc++Dn/0HfdBDJhD/teBBh2+Kq67T55/OnbOrDEPzqC7OfoAvuDLy4HKMpx
NM2B/Nq6HWZ4hvs0EbdsvhDFM8XBmKkigLSAt4+Rkoaqit921X071PjvAdse2nGKkLKJBlF4jtOv
Iw8ePRJjsoZHMBaLfpovg8UEnDrcLwJd/w7yP52XRQiWRrNLFNUNoOQo6xzbFJ+a8QF2857zRXOu
dxelipTsK3P6YDrCneoHN12uPe67zbFcme8Rb8YzUcqQaGm5rjfatJONPcHn5udzCU+KgjMipgz/
sBmMYBHvxd/WChFvnSp+yDVCCtP1kt4gkrqYuj/PoLYcWdBw89pNp+RbKbTu/d2xI6yT7V7NV164
BuwWTpdaaxNcNYHWWW+lq1nYsRJRQiJY1pHp90ytNYdXcwKXNeasVs4vMXcYP6s4iQMck0WvHMtw
WNhYVhl1i8wKbnlITXSoK/FvK2ivX+U6U5QegykEeHoxff+u0dws2Y5PVbg5/lNCs3sxnM1+gwR+
3QUhXd1phoB12HcYsDeKOvW/vBbEwN7EF53n+pavsYHIATRPQix0CUoF9aF0JSEpRdsLjQ9VzrLt
GNURX77lbi7u/3q9hbXPCoLRzaOGv8XOfcxRerEGnxgyYTx+8ESGTFJWhpEmpUNLp+CZH7Wq3MGK
Z65KtgpNybzeBJ3sureLnsHwvMYSHxoCnx6ynXiwus0zNO5emn1g+eoeobeXzTfI3xVM5jZv1ePc
7uJDpbLjgEloEv0oXC28thEqlS3WGOhM0M0xySVqnsWkZ4EMFPH9gKiKnTgwe0YhHH38ws7YGxpP
8UtILQTi2M5gwxqQzrFsYOEMtW7ENRac1pp9J3gEQQu59MwB8qOwrRLyUYa1On/4r+mlg66YMVRP
UJqFF3y2onQMcV2CWJ5Q3Qpafm7HRrYMjNOekGmnmZz8ObhqZuge3KamuPoDHe6zxc0f6UzXKa1S
yN8JQUMoaQFyEZe8wQqilSsyVlcVRtI7/IkkYqYNJNbCyXHEsT1k6RmD93T7vKxgYyHcCoLGphIG
wfpwEHFFXVUQLRplZYM5fwK5zfMPYryr0cfj8UYsxO/IpTQSjGTKXLN2mTVAEqsdWSe9jiBx9c1s
pMEf7ZyZa3yzwF7gGdWnckaAuQHUwcS5wablpie4TC5ybNdghuambSREsnaWED9aT5IrvOO4mTRX
0YxWtghhQU2miC7ux8TYh2LzKKDhe6H7EWI9okttdC3+tU8R2faIxlgsKQyLMo9Pdbvbuq2yclY9
CNJviIFfbUe0qxB4/eLsam5OAFJyU2uqqZ/0uIcM3RIYAQrdsMIhIrvtvoZAGT6ReWCgRhIGgYkC
xiZfhETHoH/rvdOWNyB6uoeC6w+x1An0EEOg24C3+U0nV7TW/EJHQLCdy1ih/KpGLIkPTICx3y6D
jtqx8a9nanX0ZuhM81eo0soODnc+2dU/pSrlgw3eDU1DgpR9Gz1HoHMfWEwfmz5ED/f3tO6s2X1V
t+W7aBYiPl+ZGlfZ37DN7Na8G0ZDMZvbkhgnTvl1W9cf4EEDNmgb602XoHw2Sr3K6Z6xvo3XrzMM
Spv1M0egEt6DQNpocTWEQjIIUr5vMsxyEX4Se9SOY239x0PrOISeqOGJ1aPNo3lqXwTGyH5/wzkl
KMMTGV5cFKWscZA/+VP7Us1nMjbouJ3NJ5F7hGK6YK/kr0dyjnQzhz76K3deJoM6uVhaFC9H8/+X
CcJzWQxtdTT3f/H0DVfTAlKr4gGWkez3HpQsoCHH9R4sNL1fn/w4d7v8NLD3iuDhsFytXlw3YYNl
xXqguhERsX5mM7gfpORL34XU7cFWOBt//DxGV3HNDz8aOScnPSvQb25TG8UjT/feQ7Pl8Ft1l1aI
ayqjc6BY80wYgDQ5lI+vOgcYVzkzAuwqaNu6BxcAYBfbTpghXfcZNEmpYtl1hbPFqQzVbYATTaAx
B5XpE5UhfC2R5cKMNYctNMaTDqn1+L47HLWydfjKWdbp6m789dJH1H7GyrzbtX9Icgr7HJgh0L9z
xZkSTP4kppR1uxOBXEjiHwzWH+lfgV54LyaPgF8om3uAfkA+I3jxYKENF1IuKyYaZEXhtTnZcnIL
s7bMro5S0AT3C5PtrAO9CpHenW5T0AQfKtyDd8FFJiwh/5jcrWzaBHWp8LpIQaFf9rwly33pKhVr
flMel837vg1A8eDGvZVfgeRymsZdgKYDaELVk+wI9dQb+TRa8ZZ9/cqeBxnOCF1f4AHyO2/13EXA
u0R7tTLo5H1vdgFtiFNhd1zP2dr6IylrfXeXDlPYQoSGihDKF4idxT7l5LuEv3NRZ3an6mPYdROX
ip55XfDShvVUhTnRww8ZyP2r0xOaqVBgB0mHtVpTMjh06Fj7y8lVaKwRJVyoJP5m+tbko0MssTnJ
aUKY6bdLDAl3m/lIF/qoRW/IoRemECRgH8CAUdQNlevFZL/Uq21NjEmTworLwHPTMZ61Uu8qXlGQ
G9ShThf57huRxTYsj4gA8X8Cw4GuuhmXgOgX3skBehitPGoCzbGLp6YGLs5G1lFG77/cpxO3y8Ce
5c1PWU5eCipU7WLvn/IS4VY4Bs3L8L13JiT1tAm5bZnj6VVqhlf3bZTxg61q8GqbNKLYo/WBibcr
UolAimSAFPz5j4ArgNy03RdWizQDv8gnq2rsEju8dC2Ejw814Hn1Hy41cc6qF8AMeeDUv+iB0r+o
PHJ9sfloQENlCNLXMYkxeqFu5wIN7d0yxamYMTsuKYxMPiXXrzN4m/7xcThv8dyZE4pddII6SA57
T20cqyrScnAG9bLpMhUVG4WRJcdA5KfR+VkZDHrGnAmIZQVjvW02s11DIYu9eK+eM9BjCvB3cEa0
ktKr62x+lO+CD7u1tzhOvRz2H4cAO+9AFdnWtz/Fl2VO+bzyTOBIZ7XQk1uAVXf1BQVxXRWUvVS0
OgHetKDSTT5TfHl1Ks+cR9h2Ue6hgjDzEMJn4lA0lUpPCRJ93VFd/eesxlIzHvgCStPyZtdQCoPs
Fku7uglZxUiUOIP2Splw8JvH/SwSylG+4m3qYtIsXiv5M4czioa+8WOuHG4KTxyG0K8Y9NXtoJE7
t/oU1w+K222MIenhofzfPpAQvgQCacwpTIiB5WFKifupSMOiNuWuH3315wWBmwfDektA0ejB/ktu
jxuMGAzAcyoVyK8vOo4cGHFwqQu48KgvGsj2EY77zD5Sh58iV6RPixc8Hx7970Nn3iuZCebQDXdO
zk1X0YiTqgLqOUuZVU46QSKEKz5yCEp1MPFKOrFUcB+Q9XJB/WVjygrV8k5R5f7j4epgx27Qtk3e
54IejIKIZa7IxFwsqUzbnl/0t96qVuJvsoEfJeZh87/hUTy1eyJTqV+0VvmDNu7EVS0w0M1E0zTe
dLRhx60f8XjcCgN3V9jrCdtDij8Du6oud7hufhhp9RrsBgtoDY2pxCvTE4dAqVa/vJS0H0m9Qatl
Als8JR98dqhYf+7k7L2w79XJld3isLbq7/hdkEv9ZPg/xoZOFEb9AQ6SJ+oPPoDQeUWAp44PIbIO
Ufct5Ozu8wb1172mDFPIJrU9/UWdxgXwweXEZB+qsTSzc3tMsWHHj/iRkeXOPQt3JlzC/obgoSpp
TxifEyHIIWO4TZivGtPdZgGsUJgq9bXF5Fab0E0ZYEdywNCmBUkqxwUdJrDimU+8AID+TxLVAHAD
Fyi6GngWgzfDdbRq14RA/mcknyqz0uhO6sHHHEXKfy4Vyoh2EKSl0RTz8Z3yffx6DDBTvc4CpHjE
8ypoFId2gJT6GquXLTsIUcgeUpDQx/kQqZ4E34183iA4AYei8wiGUPJSksDEiFIR2sEHw8LhnIof
HJK4tP7oUmzZgHBVUeFVf3/0nZWHTa8gL899MHZo471BwrO4mq8VMPoxBtaN/jnI7hq/z0FvrC8f
375pbyOXmecm3btyIJ1fpyCIDK9hMJm9FgPcIwA5P1ZhmhJtSENUFvH0Kk/fv5v42MCavUOf4ftB
mWKhwooJ6BguSe0zsfBFY/wUbJCQiGXfAnXSfqb3xbl3q3SA+/NWWrq6wbGwlJEArjeObEB7gNqS
sPFyhEYqo9O6iZ4YYr+y/4hXVs2xb2sCS2liymxFC25gfc8SbfEXhBYcgHfBuDyVouvMcQxuG0XW
SzBw77UWOU2n4XecWV3gE+Ez2mEkh9vXpdAfR25UBpSXb5AJzaT/MmvQrE3tSj5IfsGwtq1ePv8i
cXoZZ5b0M4Tz2betSbuApFX3DQSBog06GXVSeC+v5Hbj+A1vCY1XsGDOydWCRoh4yA2DxymvB1TI
FXs6UmqZJI64PEvs+L3X/3fOzivFjAOipDcywSGKK/oDSgYeytF9fEihOqgvvQOmv9kMd1GpOSc3
VeXej22t8vA88TaTmqyRsOPq7d9IHa6IIh3tStbapkQHhK4JtekwYjl93zxh3p5Be3whGnjva3rm
Pu3ulYSu9brpzXi3Zn1lhIjS6vPfhBtSUnae6nsrAMopVBGBWs43dZJNNil0aWvVzN73RkgpaVFW
e91cXEaH74oEv18PZMAyIOPBsMeFmBEdsgovzpwSZXv168j1DyDk9vp8UFfaQh5saR50ITGDoZB2
cmvyhmR7BZmMQ7lHOc7i4cbrSowimuECcN1VMOSyKN0xoIcoRVk3YmLLnWxAIDTiBHKl3QS37BMG
TDhNMjrRgCNOuqArLLjup/ueMaFskO7ugP84Yl1hG/KEMdHfkH2HaK8X5lXIDdoPrLiZQiJ8d3qa
RkYZEL7+kDk4YxF9EJv90SMztdEcxEUjE6mcLXYCHW2CU0MAA1I6Iw2lioq5Tf7iN/JkQTd8Agti
IMIKgyLXtMCs6e/97slxa6f9DRvHHVaWvsiG2PVjpaul7IfFeVC7QUY9CJsbIoUzDrsgZG+6yPnG
ZOVcgUj2ucF4j7+18dg60oyxgaoq7Frpf+5fkzmcoJYlHwtfHBH/JRByexE5t9Yt4jwF5oOODLrR
fd9V8VhaYJclVZsHxnNMBCtYdnEvdiPbnffa8w22u9PcDloudOleuK34GE2kFMkxXDdrJNlae1Q8
mHPVcPhlbgSVXcQ1zguRHT3iBJN2VEZH0TYpmTbQxnyAOlp+v8RHBa7dMcKs0FNVr2w2nz1kKPir
wuvhvgZscVfNCenI/QgSVxbDXFGQ6oKoXAsnN1aPVOUPVKlhENLlND7XQ6WzbY2JrzUYN48LDx5Y
oJQjHgcN8q6ZzUCGG5dowpWqZsusBi0RaB9I15UnQE3IruM+Efee0AzyaOnVz3Ou05Dd214zB2c9
yBQ+Vu6WkCnsRlEhcIsGerxOsvxA/t/bG++55bC1BYMB5+oHKAhHfVAtDy2elwVGgUN5AF9rkhj/
ErRLO1vTwuPFIxdETssvagnqHPM6PAixzHqlQ7g+8rtPbt5tRDNGrz2uE4q8/PPAQGueA8xev5gy
ei2/QZ3x3rd5jFKd1X2gASb63Onw9ng1q8kwxbLAg9DddZEFwb3mzasxpOCkUE9suJLkPXD+MEel
oSrulBa/BnNAMdUQiaC16dA1DegEPOrABNSjVCR4y0dVoCX2zxQBaDbtBFzvNVRdFXx6QpQOwSkY
fysvxo4Mb2pdUK1v0UqyGu0xt407/U7WDhB2n8zWNwWbp+/hvCzdsBo7UHHGWEJRmMYNZn6GxVXG
78dCOd6Kt6mJIY5rsTwnybg1nnkVvfSDzPY4/3DIvv0xsMenhfHxWF9nzyJF0edbvyPSGFlZxsJs
nrmK2W7HXPWfCNeSR910DbGlRJmpxhci1yGHcz2jXnPssuAG+Z/w+W4I+vsY8Z5roa1u4MdUYcFL
9GBDnhA/7EpL/9SHNdfulO8nd2YX3XguXRj4vJRwqm9uYr+mlaDBKUXPneyQYrHSF7WW8c6uCoyq
/r9ABuBDuKcS89h9JFToC7dsv0UOsMCQAseLvGQwRboSAbcaHlWu7KEikQzEj1oU/LVJF7btEBXz
dIV9fhtm7Gn1lROsuUMrX/V8VsusxRzjpVUqEZkdVs2hMui1opN0guOxzJ6+rhDOBHcCuodeiClZ
Jqcsqe/qxJv5qq0lKkbIKCwEyWkTC8VJoQnj26/VYUnFOhqHF24Osrwt0q4niHRbYBPc3DPdMmXW
zR15DxCM1AFznulDamyme7gtEOiOIaFt56djPysMAjucXDgKFIQI9a7kUab7q6BT8agTd4eY9j+P
WLGMlP8XmsaLIxapdGQGCI3OFOi/LaLbhZ8XounKjXW33LIvYgq7z3Hc4Xj8TBtZG35pMs3Y/ryW
mPHTAi1faSPgxu+iPn7nGherP0/+87z75x3DPll67MHRiBYByCR7iaVsMfvQBpVi7UJxb8mM+nH3
YZhygAfoHqAKFhJzNdWN0y3FAPzmPJ6Zd5fT2tZXG1EYDnUlGGkhSA2mgFJEWNosa91Zamovt/Jx
GOr23RDG9T5bFDq+WE5Vnh2cSTV/XGZEurR8NzE+Ks6VRvYLDDkTTAwFSlaqr+FcSTaGf4SDgHWv
3JLzMwHOIwmDGhI9JRebUQn8Z+R4KkiQonz6wwLA2w1KT0laSzbs2MxLr6dmv9GQEgjjSXDSGMB+
QmlPrQkcMvIm1nnOos09re7vDNoevm23rwl+H/NC7FvoO8IxGtbnd5vHR1xw9VzUB7aG93CL1pe6
UpHo9vi0zfTdCcTqYndpl9GrveYnvioYW+5hXOSNPToVv5wYgD8o6VylduPE+414iCmjI7tDPuro
E7EpS1iRTpA3rGppHDnWBcyrlq3wLT3A/4XyF66m2lt3YRq4g8Ixrz++s2fU7kKl++Z0qgykVpsj
+ql6V3AgpkBnKgcnG9EVMHFhWvMAJ99TixGu2AUW27q7erJ1accXMm/ial27P4hJddv6Ag0Vd3Kd
WF9vUcUvLmPE0SJWfhqqzyrPpIk2U+bs3z3kOKFi3/FKPPoYL6qMqHZbqxGymjIAhnLw61ei86kj
bl2Z9ARL1kVjj+oEcGr8/+7RJJ+7Ya+aZkvn5XNUtW9xVKvSrE438QQ84oC9CCNSCHREHkLA6RPE
SLE4+7xbyk5FTCDFeSlmTyXgvJ1+E70vop/8dXM3wfHYZCxV7LTBRTBRiHKa3KQbF2nhVS/hhAWZ
Wwo+4sQG6XH7bIXkokcJUQNlxH5MLzmAkg/oZZPtuQzKQbm6CJNVpW+oSU0ZpTwUeVttZIBLV1Kn
FIDBk4shCJYA5Gux6w1DyC3XWTUtx63qN/jIDg0egOzRiNZT6N7bWU8TPocGtOcrshyseY0G5wkM
G54ZWWDqnXVY3Kbnf87O9Zy2UtGm4qgEXTekhBc7r+gjNta4V9Z10643upOuEcksmy9U+1+84LXV
B2s4OfXdTq9LWb3+r5KnvsmIi1gyCeH83w7FTB3l5LwlfoHMIpq/OxA2ZgoXCsy/qwCPuw2AsISA
DjreI34kdpUUxSwNfFTkgTQMPcZlpO4mA8KYCQe54iuBxWY0NpJ7aEdItn1MmtHEVqCgVyurzKRV
ay4qAKXHPfxsRqexdbFRTgEZ241X6v3h79Z1JpRUU2cDLb9lCIMJeIZNnM8KRB8mR6lPeFsnK9oi
8FWQ2W8jeCsLAJvmImvnCyCc9QpCVZJi6BavxAU0zLmiSk4SX/eUEz5r30gfoWi6TgOvBycyfIzK
i3md75fse5MN17i1hDZDtVovSXAa1zEs9tosU7/G1nWe+6xi6if1fvKKMZM18bwK9eKtpC3KsbKn
dmg0RPUPL8Jl8eN5wzm8k3beBxaGu4HuCakwcwib283SKAujKTansPmstSGUSfAQIwZYbeoAsncA
uC7Wcu52iVSn+Fgo/RhZ2JVbPYeoikyZb6KemwhmISV0dUcHiXZTlGoFbM06Q67wP7NB7vQKWwdC
hOlcGJQUTOsJVHx5wVOFKXMULtUuRgRgdvb/1zo/GpMHrS2AvvRfLNNxoyG4j9cGyePMYtt65tNl
wfcdhJWjQP5508EmeF9CUppCheSgZ4tB7ioxpl4xtgnQ92O+Xs5QX1RU2qysuuIVnoF8wLqHkXLP
imq1ZHK8vJu0Ws+/TIM9LVBn1FDziRlT2Hy+sHg0pCm7RMlArOysYKCUViWufjpMARdwUJKJEaku
pHWTxulOKlEoelDP/kP6jwuGjxOiaA/8Hf6MO+dkAHFc/Coo/1I/m8vD7+t6SMnQ02KViibYlrus
4N8QCQ6jcdFtHbRxBVl2O4FSK1H35kj2k9L2NSCztUpzpBznHmeyU85Fui01dZkpTKVJkE6GBuy5
KVbV2jANaIHAs0mbRqVgzwaKezWf1a6blTNPTn2OukVVSmF+47DeIFxv0PojBjwtIzJLWFUJl3Ba
6SN3jtLpWzVaqw6TstHIsiTCuKI+0mJb4bH4qYOpnN7aLPzDmBeBt2SZeXX7GobG0qZw+/xlH/WH
TdxGHaTb6VnPn2kaqTPKPCTmyz0TIC7PEe8N+jEkrFQBGxTNolu1KW2mjZewTMYj0q9shlv7mZlc
g+T7XZ2jIx2w658XunjT/i6gF8G48ZNQYENcNmqyK23TSqqNC6L9j3hJdeL92DV1JDjoEjooKs8k
kzWucks9fuoi/rEAwG3emSgoUZOGy2le5c1JcBh/FFnWGyDC9F3wz7ycSz4DsZWhExen1l8gkQNl
r9MobtxH+Wp//SQ7oij5WYvVsIfIrlgrw7NFv5aaiB9+Xjp+kFJUnlSWetjPOaQX24wohktn29ls
Xfr+5crETCGKlsteArQwHqi5p+vcpd713VHYL8O99QbBi/cWp7ZdYbysFAVIKWnkROJQQSZQQleD
bhpLIw8oE6EO4mkspIx76/4nl7kkdjP8+QFEg2mcmuQ+muFwL80zvT69u4sk/i+xdp8+IYQWW1Oo
RMdGd8Eg2IfyYcIIs+clfa7LxwqGOO9LviJx+fKbv6pFbqCItXZnuv48zgUxumo/61eMvAnxmpk4
H8elDRKtYmk7zGfdHI50vKYwB3DfKXwaSsVnsBShHShnCsbYnGii3kxyl+cZquOnswfiR0ivDogh
NAg+HKnu2fwc253HBYCl4BokD9/8XTCh/yv0592kOlu1OkxgGZ0+OuoQoJH93VHhOmc49DWx8S9S
0mpktiiA92zlFQUGwuJGBizC3sGr7b2gwsBBqDPF3DTukPUu4LOKemeXqDbKf9egjzRGHKrOGh7P
wSFKQs285Gbh1iiJSbSJT2/fWo91HCcHiMIROYqDy4I6Vd21k8JuD7EKwRUpAjz3oieekNpc6mep
FKktk07zBr6bViZjwlgFSXpzcRUmWBEHMb4hiBlc7Bcu1ThiRTsEvLQBhaeTL9NWorRUmL+hvpOk
ezH6vACv6yomeCb+S3UlKf9Y3USboXSTSAbCBCSpP5Thp4tArlcXfRBccBkgPNo7/Xh1Y/+d8W7Q
OfWnl/jol+aApciElbkEN8a7XIgh77kpRoQaBpBDNJCBkqhRimCESQG0Y+0quW/zUhu7kYbtYPnT
KvOR5oLyZdaHlD5tb1zrIJ4d6MwMA+l/p2qVBN8l0j/Eazkkf3gE+q7QuGxGUVxFqqIHQwlWkURd
fo7dUqGHhUeKaPSZLv8Dy1oq94vWWebTUUF+IuyIOt8PpviRVGGyF2sYBeDim5hvSgW7HJ6szvZ7
oFciGDvLs8RMNVhTcNyvRz0Xm9NK2D/GuqpbxHVnZb1ZkhRV4YBGEP29Ro5cnrS/hUJ4sdiW3rxk
DN221aI3WeK+PEOkkgKEn3c2RpsJ3jclJ6A/wqFBN6OBBZogmNINHX0DbhOVX9MKHvgzGodWn312
U9IZTQbpxRNUwLZmnS3IPyasNUzBqPt87JgC/3fMmP4UGjVKk8gR3Z4+Yjh5Gk6G0PjZwkqIxc4n
PUDQDVXSGcg2GiHuA7cWc7OdsupZtTffiqiHsgLvdezY8XfdTSczkHF6F+cLrd3FYcEDKL5/YkGa
9gBr9jN/7oecq6WOxSlN2UomjP6jUsYUiyvOtNRr76dLs5HqqQ2y9CNuNtRm6bd599N2i0dNuQmy
y0AEWHJGC6XbT1RPxiTTRZC9y0JoDvA9nR5yih95JgdyBtY1kxRoaE6t6liWqxSBCsJ+LzyNjSm5
l+LAfqwFURWnn+FsNZTnr3tECDs1SrLvSqAW6p4CYMPFZfiKrrEuoGq9b+J3pkZr73O49UTAzjF9
U/M4MuniEg1/6CDnDd3IQLDsC1m/z7xoLrzCV0ROHeQOIGhhD18u0ryc7O3V8eBiBw51IznxANIc
ROOAe4UYOMolx+7fcR9ONeuJXBW34kMtMa2OJpkXaFd7/rHoolFwyOzih14Da+GFNuK6AJAr1730
RJ0v33c5eHspSDM0TupcRLCCXfyuVcySQEn22na41FPeWKovlBH+9AQA+exPrgXMrX4dktoH/gr2
on3Ve/R9j4yw79d0EgHmGfjTBSFBCBo1J1yubbVEExXBRm2cV8Nlqc6iDlvvOjBfORopB+Lb0BA9
d2yOI/YH1Jtswt55mUhqwHzp50bcOZ6PDC75QCvj8w4ExgU+3Z2meeLGs8gxsdWrJNx96fNQYAYo
7CgP6HLceW86ikyeCZ3eHFOeKzZYgY10QUlbynD7UVgtzVGOh2oZ48SOwWN9wJhhEw3p/+ReSmRj
AycurEeDy32xWBEkB188K3iUU9ENtU2qcvW6nGQbB8k5guHOFbb2tUGXLhqt96JjrWfjJ8cu2STs
0X8532eA2vJZdM78tmkNJM/4IOXkCrzi0eJAGePZy2rPUKz2p534HQksB/A2E15c5E7C+m61wuUR
vJTPKwmhUGIk/pGzFbdv6U6nWR53HQQtVLIzmhVwD/5icWy8dGfRE47nvXp4HNaBkcwHISRPZpkS
imMOSGhKrZx+bt8fGGdXC9IMnbySHbtcqILv7erWAN4ViM744Qo8coh74zO990jcY77kBnF4lahP
Z0+IpzolfHSU0eg3yWy0S6FhQICEWP0GVzQle1+rl5v8IN/5gWXudkoocmRhijmwffiOU7WqWtkQ
bIVNy3EIDB2dUsX9a6uwQvB9F7kclUMhkXMw3k0R5OWREzHSAtcMfk0HQrDerQvCoyxcYrdtT8Pn
L+I0IRvE5iI48HYoctlxCtUr9Rtum/PVfuEkMV9OerrXFe5Cg9I+n3qxioEsV1yh2rcOGsOl2mUA
VSW5VXYWgNlkr9usS68qrJBun9zv+ZGOtL1dPX0gjao/TSPFhZH8j70cl+1SiE4C+PiusFFeIhml
7p1ArKOybj2mJUZ70Y2J9uHmDdkehWApqp2BZwKsEdClxPeWF1VJL83j51FtZRrJInWWISKU5CFI
12kFVHtG9nuP8VSqq910eOWyQpg4eWy16gkyKRx/RSGUhEAaHWAXIEM+XKmh/I4C+lpZ3N/vrI56
akQ5trAapJohVLfC+1EjrbWQPvMWJ6EWN94jF7gKUoxeMEhczQBKN+MTK0Keq0Buha9B3pyGBsBr
1qUnEbzxtwxl9kBWc7JckblQeTaRgcc7lNYYKCQ8v0JFQSWJjco7r0XtMFI44ishGJCTHJ7ATi9/
bXhQZO9KX+95pQr1pdP38VrbCi1IJHA4p9krZ+ZkrQefhwTcYuzTdcyPzLtzY4OGQJjuGpUOxFKI
PYjI9PAH2y0cD0p4l6sIgMdkMQ0Dz0zZEZGp/XrkxdbYb0xJoDcdIAjljdMzzWBiQbdXPCtApOwR
ngC/qcFUmI7w3He49hSqfnsID/RpAcLP+5XL5wjyN9dd5BPDK4siRas+PQwzTp1HOpjrxEsSSIJ2
FNOUxErbHuSAvf7veLKQs+VMtWRlIwiJJ23Tx24Piv98H8Jwuvv5tY8lDA1W95RnQHLZOSHUzhgZ
BxSGscwD9p1jQUEs3gReC2bJ9/1D0QtzWLrtOTcSK0QomL3L7ITtERulDzF2QKOiANjM5Ty6cnfR
3QAhROkAa0B28VlSuULBQjA+9l1IS2o+ripxPgGDFB4WhOr87YWI4KeKlvt7x47FiAfNO9XojptZ
PIIiISn2wtKVJe/VjoxMKXhUPr1BVBsguUpU5eiNh+L7XaWGJu9AA8WnLsDv7j5XtG30ylyd53o7
RZtz3GRmz8V2/1daALE7wT70mCBoBnG5VsJl7KztUUBITCv7l2MTBAKaMcNBTMtcrQkAAAdIPrt0
CUcgNHjNWCedzVvlA5qFAFnXJh557DAQwvHAqyunhikYlETn1NDTCzVY5RSax5g6zatKg2JPlRJk
UqbUA6cVjPH5bEL1OGYkIoKeJG+IH9krgylvvjYFG/bmjK9rby2+1hYJUTw4wLnunvC9LuKnlxcB
P1PhDHoATF2m06C6CwWcwPy6g3Hy0FwXO1Y/91GAE+EU2cb7EZS2FtvAIuPJYpMLwDH/GoIjShnJ
FdTNDH9T3vcoPbWpBjP3bIuIkpdi+aaDwZ64bJxPtIQ39005dNpp7YmVSk4t3sG9StTzvAY6jOD/
8PW9dfLduaPmti76Ob2UJ8rzfrqpbCKW/JwO7Na/mTnRAKERI3EPg2aXv7y0inyPxj1Tml76s04X
x5bMXhl0YGoB2iBQiYze23OUOhQqjJWcGA2y1vbrxsEYdsBaNd9HULoxJ+AbjOByLtomNAuPwkAc
3/Pd/PxHYV73WPsczLgojyXxrStw+ruxBD67USZxQ1wG9/rQIDaI0o5McRkW/G9i5wY6nloXXbdl
dokXCQ4GfmiHjowTue4D+rpbxW4hoA5BFRLiy/fHjRbRf+2/PwSE8PYvpShSqW0BoOjXxayyYO1y
UHaw8oU8qvWEiqY/Sr1X993qdn+SjRRdtfHhVQ6XnjztgxqxCaNt8UidVF+7sKRMuCeudohPCWga
5b4bfsgwF9K5aD0HBCvZy1fOvIHb5UX0IgoXPIEr4033fJXiDdNyM4Rk4c66ugEtF1sIjkcJKefd
ahuPv4eDfI9HlX3UfhniOd5ygZBvbD4os5S5R7l6hllTGpDSVg6TFZMmqQ7toFnq9KaqmZHAUCLf
PgOM8rjFQv3yWkVcWMA06vmZUk1pHXCYKabKslwDZdZcsPtnIMa1inBV9HVRMuKWiEpnoNlipnqv
OvXEnrmtWKyS2AhPW1V7BWRxWD9ZjLY2+L9WxPtNGXtRXubW5H7wcEH6WMiLAHTwdVw43U3EPFNg
ZOuqriq9xO1RzeHaQW9ICNG4fTO6aJkxd9T8hd6R0S5vEg/v/k5kLAiQxbl5mwavTLYnq91K/kuV
ynKorWLsAVBzh452Bf2YugODR/OUGwfj4re949RP3wLjWdCtlINPbgqMzPwdMkrWJzvPl0t8ZAUZ
kLuI3jrzAkg6hVpO1ByTaNlPRkMCSu1cdnWR9pQ3aJghOmutcvzcLVmuqqDpBw1AlyTr2SLoUHtn
SVwmTD7sT67vUsQKUR2q47xIvF5NSzvDpHXzs3dl4hK2PLQ8lE89QFZwcBZvpCRzmWDf2otNJzLt
JuDNBycppUDSLJUQ1or0NHKGtGMc46Uchzawzc0fyWEutZ8fCz/JgO/+9FBw12SJR9goDN4kPYpo
FtzIivpB531r7d4LeUrPEtjhCNSs/qX6tTjl07fLfHmBWUQSE1nuvn0X1SIuJIpiJvq1pccIj4L0
LbtMe+MmakJz6KHqOaFnyQUoJnblcS+xD3zXLIgTpDphgXa8A+RXv0+q3Qd8rTUkC8WOwtWWR/9o
wYPBLx2C/vIRHmuwBYkCvyPnAnsjm0wPOMefAn/ykDtFL0XcpyflmPRkPMXSuut1PEl5kOg5HIdT
stmsTXc+eAvOwuIQTbW1RjyH7zPV73OPrZycJO/3O1Pg20xf5sGn94c+NoEDRPqGkmXsHuSf67+o
Pq8k3ggD8DG78K/GSX/6la7AAhkKvrEDCTDhGr2UTZRJ1S3e16LhFcROTLpvDi4OhX3FoqJesyuT
KZrhUA0emWsSzKOOEddNYQ9VhBw2Q1UvBM1Bb0eeUBd4Ob5LwyBSk55pPThgC3OtSS/Zc1ZGKmV2
4UQaxLaHJ0sccA56pfbNfQd6SdJhRniA4b+YOy0tLY9sq9GBiXmH/Bp3Ym0FyOuQM+zhNg+cmogn
TfrGap3kd6pbR2j2CHdgEgYtACelT+nhQShUKwsbqev6XyWGqpkfUO9GzPXafKGnmofaKi8/paKB
MhKBbtKJUKiZaAYGXr6VWQGpkNygspOu0EmTuKaaFIo4aGwWSyL6qh0nQqXxw9ZV1SoyyAipzver
7AOmDF5wsSvsE6YMVxJNFfSPowRJDwxmZXR3ZozesLXN/aI+4OhoJcYsFCIpSU/CTV2yAJeJnOoq
NQfoRmgMQp2Va3CuyJbVkTFNj6wZb5AfAFU//zCqIw32lf1i0V13VKQnE/8O4qZsjnArDzVibwta
4qiMz4I/iOGZsF+vFSqqwqxjyKUsB17F9D20qqgDlCZk/nYKmtPVeMfD7rpVZudIxJulxD4AWkM6
1ZkWhRgNnWxJPvMEdRaDXF9rao7wSmHPP9YXn3So6qDlhCJR14Y8W1GKZR8w6bKhZXN2i/UWWoCg
lQ81O1Pd53TdvmyOj6mAwxc6jm5M5j9Ox127/mIo51ghWt6AQ65EOFbu0KjleflOvIq1AjOUAg5v
WU79NND8rwJkc8cQYo1WH1bIojn/FNH32I3bx6DSrUPakZaaylsMNMVpAYkK5ei8NkEoBWsNONQZ
RaIS6GQZOz2uE1M5N5YWUm5RD6i1nU3bIR8DxvLWshqjjertYXgfj9ZrIByxsttsLzwCkihOrsxZ
LUvevK/GsclOQJ2wJ4QwO/795IEcJxEtnp5KuoQC2EPItSOqBtwh2MXxll/XcU7U/LI5nv6M4Id5
vfCehPXc15+MdJ5P2JvJuxowW0b1LZCw5Nq6wVlNPJE3M6Gr64unXzxowU26ejMcdWxQHROgdpZc
Ptv6ZA8HewhCLwj3oSjO5g+2VzS1OtvgE5xI0qJp5oAPbLHkgxANVR1BKX05GJJ9gYjDZqcpZOs1
RwHl9+SB1CfkW2LGajqk0mvS+qO0Ghh4Sjtf5DCgXI/Y35u+DBrHpUARvxwF4CCqX9HSvt8l4T+s
Ckg0IOz+boiOjcsKV7aEykkJJy/JYPMicWLEk+NETtEiPF227raRnX2oFNKIZR77Y+7gRN+kyMoy
7U5K3xxDDsOrTI2fjkOcITplDo0eA3EcXJ903wN14FbMRyqTsz4wHHRiDcgJOUA988yb0JVqmAnG
E1rbelP4u81FAk0uWKW69/aKWONZgOozuW+H/8VUfEq/r0c9fF+6VWMV24rc71YAdAEqYIxBuPg4
PU2dPhWp8AZ0uzi8S+u5qW86odtdtc51J3nh0ZnoYLomQQ1sjq5OLZVKbBqSCWcy8zKs21AQyO1n
TJtnqfXF5BILkTvtPmGlC+v/QfWt60oMPaPPRVwBsbVqlIVsigxFrwVovfdpzySQ0Q9cxcsbrnwV
RAN6PycAqMwEJDy8q/j08FIhFffPO/17w0eDZs2vuvXgL7gpuS3OZU9wyCXRT6zoIOPn3J0p/SnF
0q+bAU0WviFvbtkcO9YqaWD9xSAQDroLobMQ2DNUWoNRpZUNMmcwRtLPWpFdn9EXNgS+CB9HNGiw
4RVDY5Atxt12i+k/t2BVxP1C3zMqEO0pd0sKGpVoLVH/o80GmTGjQLiOdb+V5vx8fuxPqLDmstMa
pItZyENHSANCV9oo9xryFlgp0pw70WHYYXKo9yQcCJc4DIEOfTtniNdrUNoOXxkM6Pt3hG/iz74+
wAMGIn95WfVUSxKasDgBLZcqSsV5+0falNOcgZfldMAtJyio+M6m2cX1rLlR+lo+UmjkQYmPjyBt
ESY+RT8WOAJuqHFp4AxUUtesStcz+rNw0uROhnvTy4n6+B7wviMYWY4nlLMkVkeytSOWseJ+2hPc
HkO9riaE0X61WLblXFOC3bR92rhFcVng+x+Faovq50TxZuc33EZ1htdm3gLn7yXwIDQTrQskMjyt
lTplYriMlZmLHyVYfmKb/f5gtH94ysBh4RY433vHzewa1DNjNb1A3VNH6U2eNQMSIB6r0lC8H1qH
3fkxyrnPJKIZzzWbFYbK+POtJ611oA1wQeXQHov/Ce50Sb4wQ0i297tO0Bau1541PbhltwkMRYOr
tYi2Bt/lP7FPg6uUBadKEM1bTSg2V1bJ6obK/695xdvsr5WiT4/vFNljGTMWto7BFe/TPkVC4jCD
G7j9eY+LhE4myaklexIIOuBFy9LOwn9Lzhyi2U8jaYRB3V9Me2de8bPVqEBQkMiWdE6NosftpXUb
DgNNWYq1sar6wjDzBJlofQygoytzv6cXe2/YR6UezVeQ4mZRe0JN3NJgRqKNTM3TeAMpWDE3muZ5
lXY6blO7U6vh3WZAg4RBXMLNiMZwuYbxg8dDsTj+v7e4M2yaAGeMfa/4geXryFvpUMr5rGqBuiQe
ak92CRF7EkVm2IGh3HNwav5s33zXRk2hPCFlJGNwXYmnMor3uR8By1zwG5Eif+WdUtYFUVA5nmwj
jqtasWnXAGjkxH6WCrr6mMPweJ7GTako7vZf8Tu+TQ5oevFGy3DJjwQn/WVH0oV+v+4BS3Sv8Hzw
TY5WvjxFgfBFccfME6ZysgHhQlgZdfCeF2qYyS0IrzocgcnDBIhYotgCJmlc5var+Ee8xbHK+mQE
ljuKGxG93sEszZT9xH7dLq3ww2bREKmmFCnWUouK0+dcNOvnRukudpG7RwEaJjtXzE/G3Mf8NRH2
zktMNoOo15KJiXKq4bAGE9YkcfnrzaiSCV6fcKkZq9KrJXCf6QI5CkNeknwVg0177hZhlCBSUgJq
eJcvKXdsBOdnnGFeTVtmYmrPWGQD9+p9xjqD1QH1Lkj59+KFX5ndKwVPFY0+w6RvkDVQ6kRPfEKk
bEeFZvJ5punXCrUcI44YjM+A6nt2DivLZwo0UthDdOROKbKowlg480sqzUUBD8jEsFkBz9uP/yph
b4tY72xjg+Sp25AvwebvaHXwXIevMb6JURp8TzYda/RUjbyh0fzoFUFHHZpn0MRO4U+ZKLI+Yvo8
5AZnz9h9yOCuaN4Cu6qsTl2eFiD2LlrdlBjXur8igikiiPywsGSQqtsXSmIpo5Sz/9pOpIa1G0fc
mDlfVhwRkM4SNOa7ml6Mn9vB8NjKInLyXUsy57V/7IX+PmLJbZB/f1CFCHL5iJ4ZweM96xTiCK6G
HNAnvFUXmgmN/mIVMdJN2ezUBPfVI158G6VTzIcBLKMLuMy6WRoOFYjIxBJO8eEi7XRX/cu0oyhx
fi7YMXOslqNSJXnDgwTboxSa3yIwxToSfFs4DtINq+HzmzVqZQ19IQpm30xfGsXxn8eRjoxelZu1
dT3VM+NAQeyhpPHR0ve1erSwVs1aARmy6ZDAlGuOq5ldNQjRuU4yJC1IjFTc+Cxxm0hsQf4sOoe3
Ij21T2d6ldnhELWmzkwOC6tRWartQe/Cb+T7602Z4tZ8qdRCX2NFzJO7TCE/1fVbIhRcJ5gyKRc2
9JzuW0j9iDglLR8zA+XUpp4vWB2mYmecBiu5vfMJFb0LWQUBDB8u7AQKH6fmtJqW1xD/Ds7Q/FOp
AkZ6smZ6s1vmhs9epHANQL/qGXkl/7qopYp0A+kRKlGuJZ4xRP0If5u4IUUqVHriI/fiiap3zlS6
yXrbLbxF+cLmMxGL5QVsaoWQgL/YlTKjzRJEwnfAyCCyGoxpjIyZ+I0jf1/xgMDeq0bGJ7bESPPC
6sFdhlvwqmtJUSvDiSDbBY06n7R3xC8ESuVfGS3PFpvE60M5vI8crEMd8o2dpLMVEkvtEQPyq6GJ
J92tKVCsxnGzKmIBHXuJPAA95BPHTVLzQZJXDqexWS58R5M7hbX7unVJghIQK7grPmRmOqrLgh6z
XcMv3aAK0x4W2ca5zFbJup7r9gtNigFePgC321X7EO5niGW+LusGA0gAc5NF9WX40exYpHBqtubO
mHszOga/pgGxvCBZL+J5wmTROOSvJV00/7m8KPjoYp6iImL0+kfmpYs+UYl9KnZMSAbDXPPYx3x6
PpA3DXc0BQrGCqT0HnZeGXRsk/LdnPQMf5W2qhyi5gPDWetTKfd6eBMQzPH8pLOJc5xWtKduJPNL
Q66mWMQH6WjQXdE3did0hvLNS4ckWM6zY3povDvzsf++hj1yrmiT0iFhgSudlzweigBwBSbBnwXt
S0+oKNoCG8b5QtvFahgSQv1Ro8ZtQASja20YgeUYFEGyUHWy8nXpyFNAiiOWioA+Q9rY7G9ssXFh
yxxmet36/dwU3XOUQMZXEvjohcksF6hiM4c/cmTMCGHtexGmfA0u63adVEPXHDZ1vTP38GSuBhpq
mcYMfNg9p5wN7n3evnJu7elRb9KOo0ASNwV1XEoBCIynJGzuBJbDyOd3gqnodk/2p0BR4X77Bz4T
7Catlx/BWy7tZ6b0iTEOscY26T3geRZWq1+uwFk2glT7dFjNhu+SLmxo9XqV3uWwrtqgNJAQxwOS
pXKX2lk8ZHGJDGCEcLYBhO/gPKVhF587fm6gpp1s8bWVBd4nLCOU5pKSZ6RC3nSPFTtxCOUHyXZG
fcxLfHnEDERZK7WraXd685PO0AO7wn2m/ymZ0QGxGrHpl/Ahp/ACsVgcV8txsxSOf1YiKpDhc3Bb
x244XGJoJVU3EgvN/1J+5UHI1Q3OkkrfDRvxRjqCDz+DbupgGYXnalW0kmX4AVgtZve/Js238YPu
CEtVr9sF4uajjxo/+rWSzlQxfTbKS0RmJv+JkY+Jmqr5NphuRxUqJlrIplQ9hc2Cnmj8nmK09PYl
bwQYyIPsyo8pTDmR/6ET5ftWaXW5NU9QnyqcXGc8VoPGje2KmlB8rozOkdbK/ISCRAqsuGQU03w/
/2srVkZIvb6NSL8x/59mSV/aNWC1n1dxZapzqxCFBwhpDByCmcrBbZkY4tmAezTju+iULVdv7EAM
7DC97mWsWP1Ah8qxWXOMNuXApH14zPJP5H+jmL12URcVp5UqhsQ6ifpkHdzZ8jFOF9AapIi8sVRn
pGUgaaXKqI89cumJwrPphSEe1mlw7gWbdYfyFY7aq6kq8un1MB3QKbvrEs9t3PBBEUnWPOEdpOdT
G8q6UByzSnnU3UUyQJflNRBUJrNyEoCYGeEZ13U+ODIecJ0Cg84V+Wt2CuwbBpDi1HrhrAgpgDHX
mkRmadEzOCMIbtlC6dTMR5MvKz5SuBaOpGdWWjVZTmn3AyqgoIUMpR3GWSWfm8VjhQxPybWUV9qJ
MHK6uzs0C2wsupVSWc77BBtyckFtBZlmmW5fTFJhKt/axNVYzNtGOnW0SheskV4fpEPWdNmGvuQ5
r1KDzWodVuu7llzuB1Y7q+sTvxm43DY7TYd8KIRSEX7vGXVCEjugoYfQgMlfd+eZm69cK5FU4swL
lnMsspLfq5G7/i81DGdIMLnlPA8kwL3cukgNwEVGunwKqB8M7UxTP3E4+zYgcUdI89XDG2+2oPg5
6fxii4wYbszm2rRDeveBy0R5vb40nO0/gGu/ZV7NToQhGVaEPCqlL3Xw+Q9PIhtRQJ0N5XVY+Uwv
QnkcjbjXKfftDNFw/wsGtSN/YVrOb9/X1fMm+9d7scVHdEFFLMYF1aFl7Rv3Rp43a8a11opm3HIj
jHlNzt8BQAXMoSEU8/bOGGz+olNbdNCrgcj9G3FtjuXeWe5YxCFOZ1TOXpz3MSz3IY4cgDKyJGzX
4eyQoSa6sBM2joTM+lYqJeov0AiuZxyOfJ8wCsaHxMY/gih00/pQGPtoHgQFHbFAuKSx9Kb4iUaR
kG2xMO/4aY+0shjenB+Hf3HxxoYOPdkMYBqA0EswbFcWj9Nr3sJooKlVaHociD6qaLMEPBEdBGFh
OVMpAi2CgUHA1jOajggGJoBdA/nVCUnq1xgPFOJ+cJDjLworwsxuMVWsQqGk9OaV7iWfEQGeR/6L
EXI01cbX0Z67Pjvc9viYfePRbt3bersaOj61boVzWy2IZEVictr8b/rT1c1bMBs5LM89JqEzByXM
sRjPNcapW1TnNErzfDsOb4EIR4F2y2ZdfshFqdNEDZ3AKOOpbIbCnvbSGy1AwNUBjN272puQ9GR3
BIeyhMeVXaND6BLtBupZ+DZxfsdL/wYxUFoVazj0skZFMvrE/IOn59dnxOziHMaUb9m8rNAem9qx
3tM2btmer2iu16cQWA85UOII5tNCyUyU2Vfvo3kmWB4owqNNClX9o0YEB99CYX3poDTZIW21qlqX
Ja1fiGD8Kl++hXfLyWkwGLlfdZq1AshQ9U1s1vrTGfcTO0zB9qVERLtv7+m+e3Fy2TkPS+Ye38p0
n+/2VA1PknAFcb/bl8b+GScjO9EBtIswt9CqgE1TRvNPnVGMxi5435kOWeQEndKzQJaVgWVV/ZVk
CNxESD2/1aunjQpWJpFY/3K5KnIlf66zqBFRHucwVu25oyrQvOT4hkhbT9areEzA9pTI90O1ym5Z
bsP3fBy/5RvekNlABcwwiHabmfFO3FMP8yQHmRxIHt5tM0IHGpXXkLkfffs+cAA39bo4BC47gXyL
vCCS0FkqElVJ1uZjiZ+eMirRrwOp1iqjXq01sRZQNDxsGO8lVw7I1Hecvr3LvpXtBiScSPGe1WIS
2qjovvj6q91Lxy2TV0c/Gei90nF5l9fyfCEnBrjZH3JEJjLskGm5jWEe/ymR4sIZ6a9SdCvfGiLX
/Km9A4OoaF2Yg9XZsBrrx2oAoQDiwo46wsYUg+KFvqc3s9B5Iatly2Y6hOMtriIUMjJmEhU7d4TI
G8+pYst9L9QuQ1ucyIqAbhOtNZRhV6FwgT/LYVL+UpV7EqKvJxD70DpMkgrplSYFVwR5RmQrtS4B
uepa2SlmuYP2hkBTSMCRVsF2mR8KMl98VIA2OGlQyVxi94LOODUZmX+PbZ5j8WzJ50fWtohk9BCk
9vsLhrWgQ5u7y6MJUVd+YoShUTcqa1jmKcz4BXdTdTqCIMXxn352QGcPcH7EowIgqiaM31MgxH+e
RlIKY5mMkV62KrCNA0CR87WjgIPaFWOj9xBjvZqVcEJ9uFsj6gxoA1NuG41aj9/sE7K5hiH9pXID
2j6Xhqlgong7tgufNBMwbuxk6q5ld5otrFH/HGlyEiZ4AvYP02Hb+wZEiqFzY91WrZNQCJmDsD5u
lkIdHCSHU6YKjWrPyRbw2Agkh7444Ml/8lGmJYqX5DtufP5jAVJ/8HUUY5ZX5LUnsvNBLictzkUx
3gYA5SipnWUAB19gvGoSk6beqC8SYtrcB6WyGBCIoDFtzY/JDzLVvCn61MbU1dn0uMqyVwdr0Xhz
IiCFsjR/ZHeh5ajR3KyUhEm32rMNdt/W1EJqOqJTlwoaXl4m2NRHGAlR+4Ct4JKCbsC5U7AK9K1E
7Mq4Z7ezodg9VVyNVU0un0Sz/yWkjHhMCkc4+amI3yYSyh5fP++KJtUy7GEY2JBGrZy5T30L+lNB
GznkXAk4Xrz3tpFu1aRd6fJ6gPJIlcbNLzoQbY7DGZ6NPlodWsb3W8EzO41uPa+yDeCj3lOkrvCa
ZCnTqeUH8r3EnYn2Btwb52oFYLfDi3jU5EX/DULcWgoONmSBNzi2b1CbWtRfeplOJONfaDsNobZL
78s85DNo9SLogkzOpiP3IXNYXW7qzqfQjNSn/ON30StKX4o4MAAbaRvpTT7Hlhd8wFA1laDKyg3A
6foWBj2M1Hp23eZd2y7/RCwVAaGU8Qh4y578Nvpo4BX0K2SCV1G6NB0p7XO1vT2yuOOgKK7Wd02g
HEubWAWcyrE6yoawmohEQN/10ZGwN9Kyu3Bs34wHQdE+Se91lmpPKhH/Wvjpf3mo7s5dEXimZtXg
lIh3Mo9wzYRCQC6xcWLWj1ONZnpQ89Omxo67btINDD01oLnkpSqjVapM2go/kP2xPF5WUma35XTM
pAtU1Oo1B94n3Bswt+TLcbI52kQL9V01zYv3GeurgUOG1gk8EHbhesj9WcCwhEvuAFY/wrv9jhl4
lh6sl3f+J7tSivBopVTNjzDqFTKgGJlQvsTV+K484qMvOlWtWbSgHDJu2CUykNGeEAzZM0qA216X
pkHTHJGYCvM8aD6RzidQYrxpK8xPGOov424PeBZQkK0ZXRkRkc52tNOG87Z9McVaqDEwAdKJ2J4g
gpcQz4goQwiSMToXrZWrzfbWczoEC7GI2D4I96TYwrE47dfd9/B0/WRNo1L6Dxxwbba1Eu5l5b6L
2tFYSSACQpLcgmSC6I5ps+sOTk/xQyz6b6uYZ13glCzhh+n1N1OoSk0qSbitgQgl7pKzrXGuBKgg
aJfNfMWegc0DXZXaeJFIHE9t/NNOEPgPTSRx3hCQyx0Q1Dpi7XeH9EAufwz5J93388kSLXVhngiS
GAaJx5jFbkmYELsqunBatdhzc8yjWii7Lr5xNRSDb1V7zmLOMTQyufAQ3NQu8ma+4TGmmYM+Z2tH
0vwGOeaIdmmx6IFpjU3CZwGlSNY7W3wWCV5ssI8KxE69PMzX4VdBMreIBFz64ABgld9RDL1V09Xx
9e3+nmg4Xoa0msiSkUw2Ur0Cs380eys1XZmsoag4c5y+AHEM0uQpnOb4/b6R24r3gqBg9uf2EMkp
15hvxuA9J5IMdOKVrx7utKbP+9malyJ9UrxOJywrJ1xlyarPkR1thEjXu4vZOMmFJdhqJa6El3Xl
u4o3XEKkPXhu6f9ST2hwovOp8iRaZ+FeR++9PI0MoZ6dQp+BBwG167MJarXDRN85hJcgeAJxQtpD
le//zOogqNuRSeP10v4+FYH2+fJwccQZujs3SO6QYPZpH1BG+EwsFFxBv+s9NEl5EMNCNfJ8/aDj
6YJzMUBDBvRFfIw7kk+V9/jayYbCkIjv5WxfRNQapnWcXNY6HkVmJQhbj07DgOuruAIIfryZAJU4
Z8nN4gb8nUrakoECRD/WZuf5J5eGQNEEiBI9Ok+T2yt0nPLj38LXKWh/BV3M7PfzPWfLcf7jQczC
bDggCAT5dquYEnStMgBnqKSPIyHIzIk3pBqX5Pb5OfT3Jxq1bEHKh13/3dU4DhXWqbia+dc8t5x8
ajyygzEyJ8gZYFz6oebgNam6Vkk6/NhvpVrlZjYmtygrxtS5k4+JHVtW6eeSSKwtYuiLmml6SRri
QQ631o1wHruxcJGsA13qO7Z3koO95UujqAbcAC+oAj81Mk/MYGzq09CGqOlnc9j0FbymJvOB7QZ0
pL3JkVf9rBcu/M+7TMiUZCEsoBYf++dkj/Ep+yQg3kIf1XlYn+BLzQFK7VYV14+XMqkSEZjVsUXo
ro6ZWkQaagGElh3yXtLTpPNmSNLuRkdwBsdSE2sulepPc52VNvEmcuRhAeba59JaFw0NAycQTvUj
9nGM635ABlFQ8sBlEBZ8UbwwAAgxGlU3BhQDDhNIXUdb6uQT/7pyBkvUvsNFkRgIGzFEPoOCWVcx
RzZi5diUBSaf8nyjrMmfqSa/H681eWLxs+/4EcAjQUXBIRk6ajWmEOyrYe4tSwpUMIVj7oT8b6+z
x7jZjkdDBq/ISCNcCvjWHZoQGxN2U5d5ZCTkvK/bYyuTnck5gKhliD5T0NP1WrzDKkrH265KoVtV
Cf76X6bHdRJaMvwFXnuWQXUC9j4ZGHvEv6w2krBZu2FdCZnbI6dCWxuFkztmuvhuxe9bfN2XQRB0
5Pno3spOO5n13fIibyq8L731E8mdSWQl2KzDmeJ2u7Lo3IrKidaQ9RYkbMqso4F09eJfu7PxscaB
QqsMBT4X1XgG9w0uT6AH1g0vzP5ds2QgBLrvA4SXbdHGRU/YBlsTQTZJ76B6L/8ytkcqGJO6Legd
TBEP5eeaQ/wR1oz1VKA9q1J3JG1VyDZn2gu4EVHaySqV+bDylXE4JdpKc7OipocK6Lybvk4KX/QN
oqCW6smnuImL5QbSLqUwpbyx7P8QKwW0TNJHSlI7gAA0wRUMH1neTCEu5+L5frZlRNrT4z7rRJlV
XAqrs/o6ZBVdR/qeZG1zJlwl/PsBIbzqiNCzb34Hgo1vcAQbpD1dF/lB1M9n9aUDJVrCvmL8n3oa
1Iy+Z62FZVg1K1BGC8ZzJVN9LVXQd/iyBbH7FWTqYB1M/TpR0JamjceDMv/Fn2uYiFkWJnVHpWEi
i8yOWVx0SDAFoAw4b4iWlr/WXGOZNJK1cn1cy8diqRtrnk+ZAbd2ksqMZ0qlghF8THA7T9kT2yhN
duZnwyfw5zS3vv5oTJa02+JnlZFCiR1Qv9TOCC3vYk/NaFF7qZxbW6feSxVRJlhw3vN1WZkwPwcP
tssuc2pDTONkcVjwXaOKT2rqG68/M1xEs87H8UJna0HHayjx7liMzeuIbjL6mzXYo/GWMPT0YsjV
lMaV/keshabvxTXGVEyb+o6tp88sodPZZC8PPpF/Ao082Ew9NLV3LRrW88Ff9Np382zbc1ppDtuP
PlQSV0yWDYwVIqgHjDVK7BgStYJvw8xdq5nHb8VD68dS38QotVS+Bbdx5DfdZ49jxKhuUzh7w3DN
d5iND79+8S/ngCHhpkPFx77a3bgNcgh+5y+qttCMm5bffSKlQfBgR46x7XUO9FniuD2AVIKnDF/N
08910kOYBjr4xFoxh1M25pNF/BXVPlTIYlJ9sE5llgMehbOkavziRg+OWQZPuPCdJkuy06od1G2b
LfENo0wds5OFzVnYE0N8YBpRy0RBJApZ+mXHq4GlJiuFL5wHObcoElu1S1qxDa27R0XvVzQ0HzS0
12ao/2j5LPkq4hvXZ2CysXheDccRD0Q5ZiNTSh3cYvn09PaIpqKmKSufumiMzliNO99IOSz6H8y4
cHtuYik1zyoR2RTviMtdBuuDguzIHnRaXkX4AIdRwsZxub79JaADSuJgEOo3haPLbGuYUW1+2NzP
4IFf1HbjWIeQv1uO2mNXTxPY/1uyU5i6wgIUu3RXQhi97HjAt42vjB153sIN6oiZ1QblNIa4EUG1
HEiKO3+As6sUsMx/TbPalvJwsng/LZLaNWEQ0w1YTYhEZYFsNpEBVuGGQvHQiX24UEZEmaMaY+Bz
BbaMTh5rCrN/IyirSWQOwZoB/OVhgWde7/lqhadgugw2v1VIP10bZXAbfmaV6eJJCp8B4xX5IE7D
kechjI8eT3U2GiMk4+vgLEpjkmpY5VNWYdPHmpzzEGK0P77ZnEMGdtDG27tWk0Gan5Q6yQSliDdm
hsDtzC5kpjx3HGNfKh2QZ2XkA9skv+eAPKo2kDzb1R5COUoI74o9oV6hDbas0yvYS4co9OUpSw/s
rM9gttcBXNVqjE4YeemydYMyyX/WA+4C5WJVo3WwP2AdZz7RGoCXqp8hxzmHsj6Y04Vgrb54wxAy
4fJ7arirDm+FD2ljflV2ELViNy1QzomUs7/K8yi4giiA9Azk8p6YHTIt+ZlVd0V5p5qhwyOpsWSZ
2K8uC2OrJLHt32zllB4g396KzzVQGvwT+ixDsCJCUYSqSYH2g2q9LS4N9+wezbIi8eBer26WxIOL
jKtOheeoWu+wOSquPT8jeZzCMY/tKYMHH1y1hvtpL+AXLNlb9uVxDlwfK/xf//tywofEpsJuweoB
LRo4yi3myeo9hJhgrR0ckwgwPaE7cKJwWPnPdOFvaRJdOZnINBtv/BTWBEwS68iIEU1hKdkLhJaD
KHmpX95KV/F9WNELLSK1ApbH97Qv15wBESU1bkqmzTZ0+O/xwfuZguQE/n8rw2zm1EnnAd/Z2xHb
vGUyAVXvwig0I03JgF0KEunQTRwYswl4AZrVIE8pAEa3yedtjSECTXLuDExbN4IovJrUvE0XXbz6
nMrl9mQQq8Wz6ywq329rho4NC2lKxIveuzUArk9P9ITK6yhsROcDt/hR0NWNj50R4uxrFKphqvSt
aOg2nVfkLsMKzvmo5ILIkB9Xh4NsejEUibj9xAAzyD2wz0amX5rjOFr6oaCRg/9W1vztl4fR6rnu
eyEJC7FKZnpNzZmsQUZyTUBdI2hQ4VHbwUCkq+E0M4Gge+iJZrCiLxvPnfUod03JqvDaSZF8M+X0
BVTyIeitjZ7AOXzpeKSXwa9/5HX2NEsJtY46yJ+4QPgSMbcEpwnNJqWABi8GCVRpw3IQD4GMRMfN
nNyALXWvVBcaEOROKb306Xyyx4TmHMQnMaooeGVN5Aeoco/mP9E86EA4G41WXwGMRLpD6RGkKSwT
zAqaMOaSmdShjJ53f5ttIXJspI6LsP+4KOLTWpPceIY3L7voy7tDkR0gll+oA2UQKkwWnCxe4LuA
4K8W4B6QqO8iIjU9mTMmqeJFNFS5pts5Iwnr38oCcXJT9CxssA5OJSNw5fPqETV7L0+8Qrp6TovS
ajmJlEhAaEINf18LJ/5cBjhx8rR1rQmcVuDv7eBKoIojAMi9u0084xApkREGQB4rJMu56NTx2yDO
yjjv0ZvHuXf0jgRIPDjHygDLHa+WFCTEq2NIdmGK9gEf1aBhYvZ0YPQK0XAdkw4cEnMu7ASwsvZ4
f3bl9x1/OkxmpZut2aV57GyYJXJC8+p569KI8VuGLJNNSzR/ZB187m/+jmx8E5mImb23e0Xs0GVC
euQ97hP5fwgN+MXmQONa+h/0YJGb3DWc9GwAea+J+bEhcvwcLyl08RPm8rsK/Rn3/NbrCb1g8OjZ
9i1uFRgYUZTux+6339mI1xXKe7eWqtNCXrrvPusIj4IYfto2vfDsj+9+/HHqnWMDKbCYF6rwSCy6
ae2pMNTCGmd7KV1rJVFc3pqeviRBx/btpPA9YmOCtqWsp9FYL2MmMySXnY1mf4Q1haBHyxVgVQxS
Xox5J3zcIrCVk1qOlQIXVwQDjp+YGV2L/h5pxvIrL2ArTpXQOHwXvYtsOxzkvnYARc36e0fN+1L4
0Klr3u310jJ/e5/hGC4YPGXAvUQt4ApC4YrTosi8FKJ2ZlG41PbLRcsqTu5VT5VnLPEbhoa34NTF
/bkw06zv6T2c5XUobNe6GfNMDT+SjzX/NV9PYjUn0J4AOi4FFc/M5XnNYNqzg0OIlexBPEnkW6H2
Hx1LSxJfh5+f7W4QfOZ7ny1SbhNe5cnTYOLS/wxfs9Y36NlxUXUncigyjqFHfC9WoGvjwyJKTEq2
fGAXvoMinspO00rzeNa4p1Q5cTYPzgxHely6u7RsqOtKccdUDaaR//aTXpoI07qg/dAbBjmKTeGE
tORoQSaBQoMtn2w4jgbvIdG7IDSObwrPv8/e8jW1dxF09UyfAAQSyglqJ7c3C9Kgivh6RCwThFHG
aYNfaTX6BwQIkchTNRsmrfaLFqdE2YmoMM5ViyRS20meprp4jRiWtJJP2OqkMTdlmwck9g5sffEc
6F67yGms5fQPunD4taayS0cMs4+5kTv/vvkSzpBVI3GgiuzyNcvY3ymNCsyYNXc9SzPr7naVOTe4
woIr9sFQXbjGmftLzFfp+IHbJ3cETuNEYOU4GfixpI11VDg5a8I46Fcgo1+0o+lznvqbQeO9qcA/
s63XmHt+T67moW7G3jdya48ghE2ErWkNjOiLsQFgxxTF2cu+AQvDdrSp87RxYbom0QlsypG722rA
6rxZxGBA8p1k45kAVbMkD9mTueXqBnioAINFZkWG7PLkdb/5bw9rQd/OUhhhwxaoQqfc19i30F4D
OCQR3epJbibUvYVRxCkJ4KG40Xofq3N/hM+IdVFIeM3BzrluLPsgeSK6U6NRCrp37Bpb3OzjG2BQ
1dvO0bJR0fGgRrdN3OkhSdJUH+wL/Ws+T+WMPAGg/4dh7o6VLSWTq0Zjt60xmuea+a0XuKGu6YqL
bit0RUhCFmZzVvhtlImcPkCkwFHGTo6HMevRh81kr70paELjgvGjn5xFqOQGR2uwOP+kpDBQdra0
MZ/0gOrZoU6Mrk0jhWiiZkQrYwS3QD/Fcv5a4aZKmC8LVW6gW4EdfbbG8J3saYibS2+NnvMKi3hL
3qCeNORaXA+GTS3cLwr7Ulo0kkvuroANOziFovIUIkQjxaR+A+kB7Zi+xONHQNBXjd35YA/BcV1O
22BN4XwY86usIU3DmMfEO9Haf7Ixg5fHqffzxvSmm4lxLg1YMZkLjCmRMlGcugekPmaG2/gEcf83
IELjCLgRAF5/gwGTCw315WiR0wXsVhTIlrZVxVLauNUcZ1szPw0ENCinGsfxtvsAJZpSVVkp913N
qvVR+dLBToRsn1tQH3gp+7r8yjY9a7BoO4woN2mHdcbvNYGTLU93xnf8ITFb6X3K3/DPQegstPx7
jdBwIvgVzPH40abXJyEiDsDr5tjj5KvaTHZ0wveLP/Urb6yVud762JK7yuZeCTGJHGs2mL7NX6Bb
pCX22fncF/D6zGKe5t1rlEfstU/EEnXyJQ1DeAz6wdiMIkKLPi5oN+w4dPo9GHcYkYdv4yA+CYru
Kr+2Zb2RIMTIWD2j2QTIBT/nJ3Jjac2T6TwdPKFMnVHfZEAnIv/t0Qr9eUoeuPvnkJbXZgX4+hhi
wTLj9wiZyHcOZwLCAx9xiuxFmoPDxremKGVVZbwDKFwDopSWSZvTBf9WMhWJzVqfFdvLu0CWPMqn
Zl+wEQcKrX9RtnotQ5wn3oGXCgoqNvK/+9lpMtcK0bxt0DVJjBmC1NnW+aqBL1Ylsst0CNNujdwk
NGiZVlxPbP4kKe0IYWt/d3dKJX4ExN7XD4/AgG2ooL8zwvb7JlUx5/kuH1T5UYIukwrNFiTmJNCJ
+JyS7YgdXBUU461CxNBGKhRTX5IH76GmilINCof1YnREXYNu9YmoK703E6GGK5BMYTJNoof/pVqG
IZIIzduY/erNv9WGwJTqbgXXWZeMSJ/HXujNG417jIEQtYlUdPzJh5QipGAga6dxSB8xxzHmZR4f
d++3ZkfH93JBEvDtGwmmIBcsHMoLxArsC1zBtpSXKIuLP6VPza7D1PQjpn7mt9lcy2pA2aCB/FKd
AdsqhYJnAGu/DH9qinGRXLWphFdmeFP4vUKzNLTR+Tuqe5Z0b3PHfTPTCf6cxWiRjLZtuPsRe+Y2
l/WmeC7Q5i0MaZJFfclvR/8TWWk8lcxTOrGc6OgT07SXcLQtfW/1N75xz4t3BivUaV8UcO2RV3Ei
e4YeDAAbfgd9mnVwpMre3IMQPU6RfIR/prGXEqTzuq0i9fTUWolVoUzxyN3Zcn+yKXP0PkyBuqCI
+zUwuuRIYSUtKsHqz64aiKs0M41IoO0jH52U2kGY0SwKWctWG6H8biRg4vWkvY6rpM1cEvS0ueCV
ZdNIMWJ30Ca9uUm9VNFPKEtIP0drpCrQtQQSGWO9RCV/adwISSBtDc2weF6/oLX5zoMwAYZ4gFX6
49k2zvfScjyTL4FcHVcyM/1zTK3l6xUyEPrfJY0IBwK2+uvX7qmUAaiLDSW+zVSQfWk9DtYvLdwk
NkGYqLbhjit7qNzkO4z0iSi6pYJJlZP7kzM5r7NaT2I8oFCd7JDVRKB6YYxHi0zRmLDpZ1sun/D5
J3sHUA+WfOcuBVOiokydBiffKv6zYtmAOFIAYuw0QibHnODLaLHS50lpdQ3IPwUsxYp0j0ENY+7O
tk1h2HnkTKLBgojgtbrsfnUhSmDtcJPDP948jrw+RWCm4lFEu9d8hPLofhZGn/MExllnPdHRBNdB
zGGa5/p2wBEnT9W5Oc3OtYpYh01bB8//XSXjouLgIWKDwysonozy3o/eorwupCJ4TrycjvEQYFwN
5a2+AAwGEjmz6STmpOe3/Njk4CFLZKtmKAtOWEdQS0H8PzLbswVM/09TbiKEQSOBRtHaz4TY3rUs
8Udm7cWDb78hsPIeBw/IMs+2wdmIrja0LVyIa1VPLO99rQ7YGl0sQz6fkQyLKSHIZClx2BQmuGwj
AXCEQa0I3p91w1sS09batNvTSuBH283hAdAZxsx5vUWbrxpcYq9uYIY4CZ40wZBGL5J6BuTzkvC6
oF7fPHm9eA3hbC2Xd3PXY3OlHn/tj5HfVNnUdW0kmX2eg4mmsFuq2o1HKQSLOyoTYDUEbcBRbpYx
IUWTSa+tuJP6Z510LpYfT/cwmtldZQOM1MFDmnHI8i23hQbinX9DAPkfvDrQMkkTW5IcoXnycNeN
xfk03+Oa39aV+F5m/9yiLZmOEMYWjuPkbHtDx6wb92fvu5HNfMLrTDrWi3FlTOTqXrV18emij9PI
25NQMosAVPNQ/6PZO0qLa9IqMBmTn3vRbQiHMtQFQDO2vcFVrdqcW2Z4mPm7T3eZYISP/6Cc4fn+
FRyD4CrNaASW6PRmXFnAW4fC/wIuYT7eY///4EpSBTjDr82vTe4FkFgbvPRZkSSBXlkWSJG9IFbM
MkP6xVWrTkYA9C9N9D9astlNdSF2AjYtKVH0eBg+YzEI8OqHO/bTrjydu53kYq0lOOBJ2xjpBqF3
ux+W4wy2Xwfir6jbsE9mvL36lOuLPU/IoSY1h/va9bXOMQ848MbDRRC1s5hUbrYMuTPlaxxckhp9
jlW8c/ijkqcrNBGCRtzseOIKKTPmA6qD1g2eWPQ0bOrHGw0gIqe5TPFVU+cJNaerfcxeW6TM45zk
dat+Jbkur+S8QTWX1G9NUm0GQXo40wm07Ta8ektJ3DhjdCjSOc7dHvwWelaXi4XiUR3b3MYZvSKd
+dA1hSGoV0FYmbezIY4cyv5KksWYfiqkAF5uuSUS6n1BmyG2MMyFoUtPCUGe1X2WfgfyYauAqjW0
QCWW1P2GsKNmAw2V6POVXNEJSWnnco7ovlzfXXjabOYV9sf8NGFiaXFbZwMQxTEihG18lpEgdzaz
105T7zP/3VNkRwNhqg1Avva5kSpnO/c0IStiMBvqekF4b6liX5fubt//0WKOPX3WLQfhAj/+jMJ+
XUTzkXsiaMmp7EEmSulWRYroIqOtCKJwaPeUSKc1Vkka/xI0O/erUYAc0HzkMDPIMcGKGjuThH1h
+oM9txT7WKLXK1gwTJ5Mk0KNqOJiv6yhTCPQNcKCLnEcl6k14Q4TRiu65jpUe+PywtUJ9j2YgwyJ
LnfdsfGJmAOOVP+EW/VEBEFDiQMnVu5qj1yMTRRwJwttd98PzbTzWFzzajkfY/DJJ1flFBMh/reZ
eHZ/W9gIAslvIgokWldKn1+9c/UqxdKczq8b2Ya1NpmSVyZIaIp7B1zeVhYhj+Sy5kdFn6LurmJx
kdEklByZnKH8YOJYGc6AwzqG9Q0kLu6xlkFgopteUf7cdY37XkcKcLALW2rEvgEMwd+x1t08RisT
NRojX/uMR2pjeB3LbralEEzEA9rZa6R9hX8bwnPRgaQChnW8jn8snH21SYrV6fvvy42sl0GeLzF7
UyLaPus21jHMWxXe6s4EFE/L3wpb/5BCRqs4oMJt48CPM6c/pNCad2lX2dPje55uuV07X98f2Edf
g8dTSrASYAS+kqeLm9YKsjwBF/kC0gpbJr6C1xqk0sibM+D3AWjYqCoVsNVMeJ7yjPL371Zi1LoT
HrYZrNq25Fh2qdSOzVFokeU7PvjRllkfX5MX0WPPh0ywllm34szX6CMeOKsV/RFNGehuWxrtP3Po
iejyAQvRu/knLD0REpbwPttm5r9mR5xrjUf5LXxnrZ9soetdFtK19v+rQs0h1eVUy6wnvXLCOPvw
Zp4r1czuH+GOeroWoMHL9l0BJ5IvyeU0eFTvGPnxygjd5Hn7eoaHOBeV3S4jYQqZX0fZS55d/PSc
tq1hg3hz0HJDNXBKmKR2T8ZL7/m0oliAd4EyFlUdnvl847pmaYgSUWlGxD0o99jkEwcClMyQPr/1
ngrBqCv5+PZuTnGiwMbEuW868LcYeXi4oW2wst9qu3qwcZsp5EJsQUIYMA2G0wPfv4dzbxiK2Z5D
jkhyWVJNYOzfylZ6icmKt0KgKfmntryn35Va4Otpjf/Wvo60GULR/nqF5qUvnnsRSKHyJTU/2JlI
n95qYcJiBw8iRtehO2pvz2AK9DjaZ3kcbKEFfaOw3zTQWxLHnWI4F7w/QG48hvgTSGMOHNcTDDhr
3uzf5IPOF71PI9wtxsn4fSmOEE8VZHVZ3VUyL4W+7QHTx4ntxsDR1qmar7n9VfJ8kBZLgZEdSszI
Lz4VXUBRsKRI/yc+XAx1jP50BXXmAFQLQpkF7eZ+ynLU0YeDDvoiq7aZHi/yv0VGCgz+9a1Pkija
uwbxMeQxjsSdTUK4xCdJSxDuV/37hHtpSttk3ehnZliNCuMiGVhysi1akJvsHXMxQtVy0jG5IkCx
4lq3zwmvKz28upFMgKSfmiNbhufw/bnQFni0ay0YnFPiGch5bm/cHeKyX0IxlQ7gR4dGyuf82BNu
hBTu6bxuSGG/L2h2pTnHG+SSrqKlrywC3E8w56KCJUZuKzcdRd0sSgUfeq+3VT6ZrmS68Cz8wdrL
KQuTanYPTHULkLGfVTYV6X5bWqT7SabAaWmqgQykfPkjpUmj6QPqYZSEKrH/ZSzptBNkwXQaBg3U
sW0Df8HoMSaOeIeM5vPcOGJhXezZapv6JX0m+025MZDRwSQ1TKd8d67GTvB+Vg8R/+5k3e+uPycv
O77bEy5Rfz+ORDPNrxn2ec9F2lGtUXjqXNnudQ6VcNx8oSKBVZS1po+6rhGpBDbyvShatGaNMc9m
CcbySivncv6hE9ffSzJvPVyv8dLmIbhcitCM1S/a0/8fwU+gY7WaRiy0TGlRXDXrP76TsihdcU97
uKMcVunteceQqX4AqLQyQPH2wQYQAZ1Z41dmSeL/92Nzy/SMExFZJk6gSqqMC0S5fKJEVtx49JsU
bmby1AoCwq+LzR7EBSwv7ygvjlolHLIqwbdwDJoeNTyf+3ISCc6g7TJNxThaEtFUKxIp/JXMe6hZ
fFFe5sLARRgJ+yHRT3PtUBiBYXFxS2r/ryEMCNTbfQ491ZTcynGY0Yzg4r7gh4lQCIdzmvrHxKDn
wYI7lk6TI6ZlQguC2DHpivSJ5Y3XxQrXZcHjKK7tPuQJUg/mslrcaE7H5ASC9W1gH9QVbjE14NT6
9HJVH0g3Ei5owgKefrrqYPkd5L7rPRpG46mgBp2gBGiMcCNkCdrHy7Ka6SqpxSbN1XVJ3pfwuD/t
0oCRwAxC8OjfdyysJzZq3dGOLwyWcl5W55RTEi9BHHq66G2+8UlTlaC3VqYlIaheKium/2xlThPi
EoQb1s87E9+xQtbugMD73Ebk7vEYolhALb8ab/jTCo11RDHswss+nnKoz74X00RJnzD1+omqR3Hg
9G90Cs4pAB57dPVrpoqwR7/HTwO6jXZe2Gzo1/iP8kSqi7sEILnDqqjRtTPMWFRhXkXueiZRKs/p
E1jXJ882O2X8bo/tHQfut7hxM2ARERjlCBgUORk2uju012+y5Vl8uEOiRYx4YsO2kGZdD0hpeUyM
31Cw4TbnKHM+mKfe0+9CVRclpfhmaCVySscb4UFglf4k2ieXuy/Iy06hMxebkxb1O7cyDvrc5SMF
3jNPehwzThD4nKOxwm7N960HSuwnEIQv/6j76YE/HSSpxVg/mlcae3W0lgr2MPeb6l37osfEj6KT
OdpbLwMZ6Xxwwe4oM5GB876KHQjEvNd6A9FD9Hi2diTME1u5BDdHhmH+8O65pDJcDfUG4SyxuEBn
3K8bC9yJ6WLtPoJKgQkRhqEf9LionGgRjESE8wWuOewpCt0xpHlhZgpFhnQLL+V43tulwWERqO6g
qISQt4QDCn+IuJgBWy/3s7q6WctM5pF8JfX3fd7xeKT7Kka9/jy+XhzcC4C2UC0+LoMgFJha7iwY
oziiZykIG6KD+zhLLfvNA+gIL5nBb2kMPwaQX8qNXGQWJt7ZmatxbLUoZTUBoRUdKDjV0gfjZWVX
MKcL9vN1uwCi5b2eL/PBp3EI6Jjcb8ZtVuZUgyjvWt6tOBklmRemGH4NSoMm0D2iOqXKjbKCrFIh
2Dloqij58KwBOESi7xeN7p1jZ+ZNLdcXdCYb52pNRgJyyuU0jf7UvQKU9obTzi8ZFQVoha1leXYT
kC9Gb/8Ow2FEKwXQBYG6whFIIEQcgXBfO08h5FcUKaZHzHJvoSnIpg4AupKK1l9yPcUcTIZCYw+n
vdA23UaNw3Unqv5yHIGNY08pnf6XQ/q2GK3KtmtkjfNArsHeVIXksSmmmIlF1+SUPeCbLWalYka2
t7lsUgpCLBGXblLkAy+3bH/k4ufA7dkMih15kTo9+9ZmVyPeWds0lmVVBNfOPd4IVc82SyLSmsZW
OlDs0s3FHwxFa5YoTZLOyzuL4/1exsHMwsyUj+UObETjl8WxR2ojzTphFYhXWEiRxXfVkE211Eo6
6C9FPK/hTE3nptJbIiA4TvQ1vrhRoaTIS/IguTDvqSsoP2AbLBpAxfWg50qaLfLYeV0m2qOvNu5C
SmjWUS9CT9034vHpBvAF3A8AlXhXRZ2pXCHLVZ8dTSncxKuaFdHnk2ziBe7zy9SibEswF/uzSk/n
16yAcrdqd+Hr1AqXksO2lx6LANqaU/smUkNzMO4SSGs7xvUeKCx0IbkYPA07jxGuqj4kLLsfxQK5
6ybhAZA8igQ7z/NdNonF/9gy1eCyO2cKelAw5Y+qk2mk+Y8o9BCgkuffy5nSKJTiZpAlDXTbgqGB
xXcRsvkKN/HxiZJyjNv+7xyI8/MH1Nlzpjt+spTY7Yf1yymo6A8EqoSqlqv4IFhI+fd8dWgJc9jC
BEZsUo0EoqVCCcpEir0+t0eqLeLojDXdWd2mf9IRbvr4h/vWu2Q74gGe0zgutdTAFMYQEcTQxSVJ
+dZ/F17v1EHb2QA9/XpeeZt6MpIxfCzXO964XZR8zbjfCd8tgB99m+Z/eA+0UuVTAmxdelkllpWb
6Hpdlu8hyyL49vlTPZIsD4n6x1vNgkpmLtqBm8CTOWH1LesSTDx6ekW13QHfPrFv48H42lo8h1wT
3ldunbyFHPD1Mw+TX7MWsPkslgPzK+/95Skl68b1hijK0qBonFa5NPTifu8+J3vyn/3tP9DAf89N
qhvAYfmBpLcqHb3eTrzREugTMZCsEOXb8VxpirNDTJFCEHV0x9Q/n3u7ehh8oLzgpZxaos4Q+8Dt
554erc5ucPPJsjn8xlqMnQUqBzXV6OCyERf9GUw7MjNqnLFHSPyuw0Vb1kCh+sAyZwYjlwzzUTDk
kZcQXdnS7j0s2zssMvvO6PZutr+nJuiseTSkhaYdoNj30DhYq0/Yyfgb9swIRsSq1sG5olVkD/p9
iLFNGe1h5WljV8ZiAFKfE44FyHIr00EAkHoMyKGHSl2D81mkIhnx9XPVJjcE0dyMGn4w8H0VaN7o
TOi+dPPr490IBStmh6fNl+MA84xASSEEfUbdb2F+TX/VBYct4f0gzb9JTq3EYYmioI7jYF9lSX/m
hfh490Z+nCnFSBAC4h2XL/Op5qVaysKDUxQnGxbePMhixV+CNu/2qQOrGWf5mHkwjSB2U1GB3epG
5LiytzkHpiwioZlzJdkciu+1DFSOMy4W552KH1lIT3QrIAXrakR15Y7PwTm5Evjsz5o2GTgAB5KP
jS3qECx/4NfL7GxafOVHVK6fttJMaWk1O354KppuO1FzNT2cpscafLGojPQ4hOZy/ivnlVxnMkZN
vvng0LeBhxCN0YyFprII6+DdKReXxOukPevHaUYICZpZaIxnTUzy+XCCBwl/lKIydyDf7DKyLNR0
brcud8HtANyrwmtmGxDubAiBJcrMssNmi6wOXOgae+CiuVp6yzMMEhgRmMBh7GLMZfVwGxbKqWJR
Ek6qkCteHfH1j1TfreLRvXWNMf40HSGkpY75wQFE08+rUveaLF+yHh1qo3rPdrnWoyAp1GkrrreC
05t4ZUMoMK1V4CNien9y/XDBI0Rklf25B/xdP+CiWpG6vApsnHhJ7ZQKUQTrsP20RendvRJIF44d
DuzKT+PS3W/k67fCsGMmRMbWy/cbkTM/WkW68xD3tVEThSYvGHIpJxpdvbsc+Iqc1Ah5FQkJORKv
0HbIvRMR5S4LrerOSuPA5C/nLN+8KgIScY1bZ9pY2YUnvtgMOxoRLNcZgOmFnWN1zJNm22cJATjQ
ZxpcgMLgwEekuZB1Q82dxLN6UoC+F67TOpK8vivcxxvGkxWl1QJ9VqknwKEdI0zR6pGkMS2eiknu
K4CnQV8JjsCwn1tg14AiBWF1Txs52nP6ZoiN0ddqwYzjOI+z7L5v6ylQphF44gF6hUPngIad0dmX
6gWXuAW4D6maGiDbjRQsDtcDwLNJXlVGp58ajHYAMXoqGPvOCkziC4pCbfqAOHsnka0jGWHvABOH
PLiQ9OaALkXkKxC6UOJfFDWofgZ1GG6kbb/mX7TT+oLZ7IIQhYgPd7te9GvkEBDfxh99HB0TuNnw
UGuyvXYh0cZITtAGv5SPXXmX3TsxpfkP+XS8HWr+u6AoMHAWpVrXL+MY1fTnl835H98qtDCOoWXc
ch51ZQ08znwAZbOETgOiFQuUKzM1MK532BiMq35ZviUQCJuegEZvK40comtEYGQx8LsmjD392Eat
JomdbypECZ8G40V7aZSLEzr+0HN6haFR0nySR4T6hEoq8x5Bm/jQyGf14CxEtb+P5dWIlWRd+RJe
EaDhD+K3vUUSEi8AlOmOzY04PZ/E2OS9GCCygbTZsUs4rBER+2I7PqbaLFYXO6ZEF2xgtXY0n6LI
LH7tPbisKl3K70F9vI5so6WloJwzY1+W9JyR7K03QAPZ619kxe3OTJlnvk0v2JsLdoYFjqMg0gqF
nGaWLRQQh3qiZh1TMbnrn0gCYclD9l8muyJp9LtgjeRw3kCRSX+g8VbJFB7h6j8KVDR6OOtBcNdo
YVa9AUBet8fUnBPR4PNsxFR0bIZK+rM0QnmY3VLUZTUaCG/7YlnblZkSxl2qzn6riOa52JecXTMv
q7j6pbQleJlMt2nhUvIWezsr4e1S/ND2Drkm2yiDBJb9B8bn1/jgLZSFgLz3lJdZ8lqYNEuwXGfm
NDLrT9CAvN15Z7YCZ6xRKL1o4V4h/dCVS6suGI72KezW/8tApUISkYDTb5qTSoDr4YFKbQtnJCVw
CqKmbYnqAisp6VOyw4iVF36UYm7FM3U3whGGg60LvBTArpmUPx23+djiYup7UaBm7ifoW64ZRsyp
Jk8pKHGb8cto4v4T3ErIgrBpRi7fCpqYSyMkGv61LFcIn6K78CfZaS/LHIGs5NUrNud5zNzrgTeU
baqmQwMpwy7O0SKhR33Su8HS28FuDcJY/szG7caR8hE8magO3QS0kBGlcb0y+I3Ru8fLsmX94F/z
JpzgoHmqIHkHqd6OyUOsQl/RROAPMT6wB1Wn0HVsUv1OsFrdFjYrfycbnQoopgoYUHxRLYOwGsnc
LaaWbphdWq3A2LDiw0CNI9UUgh41MFWZx0nb4W4iGzf3DxFy4ocduD0R3xl9uJwhOa4BlrV2OreC
7nZXdT7i1Vr8SgrJs2wX+HciNkywYVE7vl28mWtZT3nIxZuRgDht/kPbEgTk2ZSnJ9Q9qSEoHG7E
5Rj2P1pdjGFWC4sQqxP+UBo8voYR9zynmokrgyDDgXI7/Nj/X6jNN2wDyDX+K/vv9I4vA91cLVPj
bggPV72HrU0kTJ+qnncj+BkSCnzFdmhg8SqbW1A3TwHCmQ0lCHkwRjdfw8ZKB5A7uLdw8wQLa2Bl
jtcc4OBbJ4jHGjp8eNJ6Ron6whfxILTBlsquLwhpny2Kv1qKlB0+yI/CEwf/alJ/wDKQphaeRJBv
hq11RJF6qp9JG9Siah96w4mVI53PSmbpLy/t3a+cp8WkZKo0SM3FFQMJwYJ+kJLTZwcJ1rR/mkSe
YMftP47eNGiGisTbxdscjplpAx4c7x5o1Ol1haqkH1lP70vwUsJOVTHxNaVDKbuVz7GBwKKW1HyK
4Zp8+APLiiPEOsPLA5/tusUxW/4nDxxAK6bH914moPLccp+GCYO8xN1eKBQE/UQn9mFXk+SVZoxh
2byBmNwKN+QAIyVjmEue+iAvAJTUtaW/ZLzfrPyf+EVLrNAjFpKHhrY4+pnD3846X0XOUAbk0pFg
DImVcoSdO2B09VbC8J4+/xJ6nl2zwz6ec7YUdJGwSWl/ecz77rGXUNRvmxFCiSS75Mq8GA4NI6Uk
1/voXW0dpdsxwRs868QG1qohwqFv9QbDxUDim2GGPHUF+rzU0ha06+tt3ySViCQWjYytpJYFJ0yz
hai4c0+/D2JfYEi/9mNsJJcw+WE96DtonC8KdFbsUyl/B7mvVJuHLfdG2BADcveJKWNoRG/9MENa
7PLSRBCVtfn0VZAcjO+U3Z3fC41lXPHFhTsXNj22u+cQ4o7Y+dvIAW2lz5VqQyGxtHE3z6YZmX4X
r7ZWuRsqBHgzqT1aouzI7X2EFkx5ND8yAmk7iIUXcXISClsV6ssaDrI4vqNdf79l1s2kCcSa9YI8
xfQ+kumBqluU7WOwx3aWMnzKtNRsIzRNV9vUb1kHDdrA489mRIREoi4Cs41p/P2CImaV1Sp6W/uj
wSxWdM7hlN/3fp108Svqpzh7REx4Je76Quxr4MNHXokHXpyxDG9+I9DKWf30I58s09+cSTbbXBC5
nOG3e+c5SW0LwxdcDd8WAhK5NnQgwArAIcOkWEmADlNkpWc2zZm5z61sGluwbRdlPdIp+DVuVGac
TXTfI7QZ4PnlUKVpQXL9KI8Uuf3VjMDfExKaRsC8eebPxtgBIgeH4kyEE05wx2BR66qcD+bUTTRF
rcAJpXqqnchnYf2QQV95T67R4PnvuhuJd9qgF+X0NhMIhcYInXfNl4QVvB7KBtX1b20c9ds2YX2h
vL/FvpB7rHS7rabiAFpJFr1t8fPfZ2AW48k1+j4xPfvLka3hIcQD4dFGOzTriRyhjmMP0e/wV61+
LSBZsDSLQxs9p0bmt25yW69kYZXMB/bQWC9RW4OON6gmzO0wliWG9o1axX2r+OBfGe3b56GJ7NLy
Q98PwxdgLZiiMOlWUgYMBvzGuW+/6083UmOWp5m0gDQiHDIhu1c7UtL9R6e7w3MmLWwAA+PAH5uP
Dx9AdAyTsdKg83whmh6VWKVwMXbIctX0yHElc9i9uXsQ4y0200QH98UfYZD2mpnUt1mGJw3O0m4L
7cBrCESBm50Q6vRidBWbzfg6WLg1gd69r9xBiQiuMRh/Rl12C4zGk/FirOsRBk2YgxbLwcc0Gy2j
laxHwiO5CcXZpu0pcUe7Otu5TqYWvYxfPnCZtCHPJroUF9mhtdRuPcg01f2YuAqQzAf2n4A5vvDC
X/1UtRsK5rMaxSop5CQu2lmnVu05kTFiW7CVvE0IOXKsDg7x3jcH6LGOjEcduHp0LFXtVKJ4pC58
dyVoWtkXQ/VS1UdgA5Yvr4z/ipprkQ/3YhAP0ONvl36nYPpgcG8DiEzOAJhHM3033wYNMRXuiIRS
z7E6MWm6+n2Jea7n43hL9XG1iQ1BYNANLJGOm+gkJhlV1h+PWS9ehhcxaarAI+2O0uVhcpvtCJ1y
qOVX0ZcCsF4yaN5BeqxtysLvS6xV/+RlXY5EhZ7NYgIjrZ00oSqXGXj0QMMG+CpWTTxPyF+14nVx
A8nF76Efo2VbLeyRgyrl/gALiqiY7TjLH6tZYYi/Y/ejfB8FDGI5f0r8yDKTWtKfj83cCBa/k688
Hg9SR11g8Jpq8lqzNFD05RQm/WLlJ8Hf4KDMPdKM015E15ngFfQqtqMTnyLWC3uuC2X7DzTEL8fE
HP2dNuBLF1VHCOeBCxIeAbSI0wqFRquaiaNOP4bi0FfdsfHUC9W9CRTk7TZKWOpm7KefPQ0kk1sv
E6UV6lGCkKahWMNYp0u+bS3YW+CbYPnB/YS7ifAyLhHZ13TEYh9Afk41S0MuvVtRbjya4XIPEvR2
IIl9IRXgcoaKNz2CtWj23NAbJ8i/Azhsq2Rw5vHL5BAiyHDEcF/2kKsQ3fIXu/ZtwuOLkI6l7hvk
CaimrjO6LCAtAMcYdaYVrRILgYNFuTirWOWDSKR8Xo5GbgtCnDBgJRniyktyFfGxtIzPU2JiQEt3
OsL5NIzQu0oon6xPmTVOyeVNK5npAASeY8DZ7nGzjUtDnN6/UnmZ6cApB6OaAirYGtpbQMd98XFf
nGjkAeU0VDuvYt4biy8HWW9+fJY9j+9nuC2xXeaL9cJ+kJwDarYMIDQRaBw76i1NEwdeqcALlsvJ
2CMUBZ3OmrpfWbQG+6PPhoEg6Em/NxlfNh6KCswj+NPSmljnQPl3Siv40lN/MYj5OWJlqwy9gUeW
FqzkGy9HbkxqeGwEvgDqegmVGXGMpYDIcDo+5fPCLdV8poIpeuH8hK2GyogDj2/R3+z7d6DQSTxk
Xb7mhht0BqPc55klWJ9ndiWvuvBaPQKgQzWREg1v2crTvSLy4YyP+NAgc9Sl2EQta8FFTWcAw/IL
am8bbQVk3jczN2duB69SnDz38aa+p2zZ8+yIurKAXXUPkRWpxArO3t1RSKl4X6PazU1cocnBg0lf
ervim+Aeq6K41bTtzOz28xjJmih09UoNTcr8XVClsjAau/+QRl1GSfMi/IdY6/yDgKQHjRe1XKEL
DVTp6trnwaAO4LhoaNUqir3BsNfst2RsDdgagaBdQfvvKAkOZGn//NqvCgopvN6l/Z6ocEUmXXoR
mCpusmx2iHP645XIcfLD2so+sAdVieTkaqKvnjCpphP0S3DSE5Y0kAyI7uK1hh17buzFzmAYZY9t
no/bB528WN7rlWRio3QB5icj7Aabr95bwbxNPqnJubbXaCCBu8VQTYmv2hLbKi8ViGCtMkpgym83
RPFluwfU0Tm3gcH7YFFIXE8wAbb+TDHu2CwUWOdMrxgjmeH/WWMRm4ppJKjDoS8D7ca5IkZCtI6f
ZYzw3+OWo1rd+VD8Md4PmGXRmbWH1LqzT62+9Xm0yjpB9IF4k/Ck3O8AzrM7Hatetke3f1vKE5t5
+NsNjZ9iRv2YFinD+4Tuc0Nf7+/HYRUEQ9I5YRsjvjokK4kf6kOIKGzrKJzVkQCm30eZsjikGdlH
cmpMaYPmO5oRpTzQWDDhR/P1PlfQyGW+Wq8utuobG2UD4263896AFBA1ExrDXitaivsC9Vd7Amj4
sVLA/1VYyubv6hWALtx2u68K0KtW1RXeOZJfOhIVr7yV+4Ah/8H4/TAs1FX6SE1dFZaT2B8AMsFe
58akAW5VOj7XtTVLULocpyFgAw+ys5NyxMx8b02ZC/tHrXbDNJej3UIPzx6GeP6xIkXh8pqy6Ncu
s2GjGDg+8qTUlTyrH2y9s9gueE2DUNvXMmq6cTUE5BqQd6rqqdZYFWPdcENYdTRBKrpNljutvp5N
zAzD8l2+CJBxoaOaIYOmeCJItORMbsPttkE6SU2zU6pkKSJD24DTrARew6al+PNaniU5Gc5LKNjN
/EhmYPQJv07QrnLmFU6F9TwJHMrkKXWn0fYViGXdVBdj7PSsp4qBs3SY/2FLuVn6tH8J6XxY6ltV
DgcaXCOy98HI4i/SrcwWHRM4AcSRIvhiJHbYKAJpNWTOd6U+t9Wt7RqTsQkC+VVeRCnLib97wHHp
to0oPe3Ka/Opc7R3ui8BoBa6hJRH3DBTLRP1MMP+yAhuO4/sLuU4sanU7SpkZ9q6zpHehs/1v6jL
19oE6IZo3Hj1ObAT/aWzZ/6tSVHKps8Qo6lvV6F/In8QI3tB6qssiMlNSAKDFQ8Fa1yrjXYtA3sD
zUP2+TCD8p+4kORJJTDmpwB+IRQdo0Xeq/o5bBAwcPffymB0mxraWLgtLYIdlwN/BHS6/h2bFJny
z8VIl/V1ePI2VAkrmfsk7tz7pu/GCB5xTLjpZEPsTWIgzeRR5ZHWfBTnbyTb6Fm504ZEY3jzgewq
gaGtKbBEapONqd7CuYlyVIsL6BQz2EtJdnSKQhddzIy6QOlB4F5ckpIyhhOWWQHG92essNEHh0PX
6hit1QgQ30M1PzlnvyS5jyde4FoXjc7d/bweUklBZcg7/6GiZTgFnChjPakZrSjql4rwDrpT/08B
jfNiqCor1uSvrxyfS+aLR68ydnQockL1EDHaF0y8D2FxO/1OjHp359fvEkjvJFc1xjOG9Qpo+R4a
M8jxYDUVpIjK4J6kzH8UEn8WBTgrtrMJXDm+PrvWZgd/aww2eGckPxnpLm9+bRkbC3y6qwvDsPm6
rKTgYWLZhCNjFnMtbWRzZUhrdRPq10dL1WUTXRbgrYQIg7JLzN457dagRhv5VGVTU6eZLO8ACpTX
ZLYv+f7auuTI+R/2ykNdHvlwU0mM1lbGlaB54mUYr/SqZ6/AwOxQUAl53UohFMANCvBCVu1Di4a4
UBW5RFT3NubOKOAK+CZaBwhJA+UfPjWnPugb7QUfdOkM45feDyO4mudNqcO+PxDicZvl+yuzfLot
nyBqGvDOsGPnBvyQ+3cdYtpoCy3jxX/uVxSln9gRU8/cHmGotPOd3JFQx9aWl+v2edlJfWJ6B21z
rxZlmpTk4tlR615rG3hWcNWPtH45OGe58H9foeCdNAK8Dp4jYguvkcEyRqSS6/0gW+/OxUXvZfbV
heq+W1DIukOEozDEJTlG2dBFsZUdKgKjgiWUVDGeZzag6Ie21yw6U273vQRnAjmsymSeptycUS+6
aKVSa8Ynu8t7lKuJ47XJo1a43oFp+MEL301YSgZtLvn+V3UDlbqplBMCRpVkL/ylq7336aPPy9GG
UkoNifVV4MYAi1WQqL8k/CV3K+BOXA9Wpnpid2kq9iK7gAxZo6ep5CJZe8o4mzA/KjLXqQ8Hg9O7
KlSjC7CapCSJiwDu6SsjPq7NxwRUB/B+hoYTpZeSDewzVcA8jUn+3E3gn9wo9mitMUMv7k6SuhGA
hkeq+c5iNGQNIuIVIFSg+kPN2odHhTEMru2JwieCF66LROEQVHE4jLCmwgqjkIHphkVOJaSz1HFb
CPvV7A+U9Lr+0scdCCxbOit11kj+DZGzDCHhRVO/XAIdjeUN9fcE1o70SoDZdJn5mPffzdNQKQtT
TRxfJtgxmBtGHkR3mEnXE+/4ztnGF4lB9opO6KXudnHtqKO+p9NHijbYPczKsfayih4yL7gX9EPI
vfe5FlT/PoF5+A4RG1N/+RIu+BsktpDITiDMYdzckke+1N04saxcUeLlLQFVmy/ZTmdPbPXheUkA
ovSodInUFfAUlVcR2Un/g0HBHVYh6qgNiUNshLUjQIT5eXbSDypTwWPqrrzzR7pfZhqVYkcaFJ7e
saSp4AWqMRO9fD/R/K2Oke//b1AVkDzrYSIs0p7PlkFZ17thi4dZH5ZeZWk1Bm7XXTx4IfdaUnOt
J7rtbQd916crcZ/BrOpkymE85gEY2ZSUYey4kEm4ZX1qClK83zLe6KUHtodAbu7f3PPZLFXfvjAJ
1gU7YdVMV1zUaEJFRxX2tyyzRpuWHBMESmGo+CcOy+AnnzDoHYJmdAqTeQMWuiZwUYT36uNex9lP
tA+ODTbKQYoQ3Po3PJwOeqseZwjQvlecUO2C7nIddl+a899fHvR2gURd5v6gUvnTsxroq8lGuqjA
FJ9HkF7lQmh78oMWvbpwfYBeKF7ITSaH8ZVRTvCULV0XbRJTnsZyAXo55l5EhefGMPWqXLq+wIMH
yCPJlJroCPqPogs4UGYarHiPScBeCmGFlHZKE5loB174ygEQu0bCxMdD4a5PVXgOA46vQxoyuBZ5
MPJZrQ7ag1V6mN1O8Ho/2fhOyxEIk3Ryhzr/ucM3bYvKNpTl9mTnfQAglFLlA0GYvIZjXzBtSipB
aVm0wZBHTkmtYRaALtJospStdLZt1nHKnNUrMVXK1p4Ou3a7nIzIduVo8pQlYEKbLOajLVEm4j6k
tWjbl6Wq3baeNVSUtXEaJ5+uNZGJRTuTJ7oRA+dxl4fqhproDs/MUP4GnPizLeXg+nbOTNr7m1lU
p4gWyQ3ZpH18NBeGCtPyZaYJM1jy9QLAnIIkiniVK5d2A08OQN1Ezwj6fhT5IYWJ/sz+k+7/d7ev
M7y7lB8oml7kIMv7MgQTTifpI3k+xaAiWlCL3yiS+B3d77IyW/E8sG3jW6LDCnYtX3ug/qgeY7Uz
H6jzAfxXH6LsfLA64hdCTosBv5vyblBxb1C6YlD30YXe5K1FAOLogzlFRR0WYnpWK9LclyQXEeNd
q4xTXzqVGYFhVD2v6lCC00A6jJveQr+FeM/Jfysiuekr+BjqHTy7x2FZsMNDCF5BPf/dQVVpXNTN
gKzA4hWBnqd7vWlzKOsMjASl7fK5oTAGi2XEUHsToRSz3ISSvXDjNv5BTRtNCHpOzqzmPQoAvrrl
0doacpQHkwaaDtPlGHw35sqOU7SpuQ3V0ma1O4ORZGrsFDeXxUHCL6TT9ItrgkfERkWDbJIbTJRD
BSL/pe+6tyt5GpkxWkbZgny6sGkRbVWywdqD71ms5FbWkDPncHAdLweENMxmOxrdptFxHdZzkYXf
7YGIsIZqH1omzj5ozb+YN36mvV3yefvjva0pilggJfglYYosXL4XjE9gnNFFcvk+qXbI9p5s8Peo
BwZAr/jL2J2CCKGGq+E9Sxl1eSQayMAzcR65thioSIChNRPtureIe8BCADqfREFfb7pPXwzOkaQl
iXP8MLuJ4YBGpB8fasKKuOQ4lRRqiHgO0TI98BuS20RSxwO9u3TPWcFxKbQPbDLGKMZEbpLZkcrq
2tVpmpPscaguMkcfwSIMIAUkL3GzQuZHlRr7gPfahHXS1SN/7npTErwXjNI/eP7xRRtr8kQA7URW
akdXymuTE7mHvvK8/b5+Xf6aZ5Ty5Pv774WNaxX9m8PzINT4IwUGR8wZedPPkKDremwpK7duyS3W
gsi6TNM7H+BWugF9i2L5UO0gLMuxK4lkDWNfuYywGFTIl36we/MNEkXpjKe/rOWqsQXyLlAjKU6e
GBCiYvQKDjGMpoRlCmSdYjNVf4/Z3XCosx2c4vELhcqKbmjmd9hijNG9PqjjZB6ziSf5GZtUaLFa
vFv43TAb+qMU9fUbDJNRJSD+Y3HhCRXgZLyknDxreXWUrZ4G0C76yMBDKoFR++9D0umvt08R4KN3
cnzfQx/O14697o4RD97VcYHiV/w4czeqoNFpKgzoFHBX2LI9YpnKlubUxZyEFK7uq+ADCAdZUUcL
mY3y36lWJmcPY+r9NBTpNEIjOux2yAq3KcJvffNfNlyUaQT6+Bb1vf3MN0FTCBZ0pu3Oa0PpWBBq
tjFSeWQqUFtyoZom8yVakI0eIjeYh0wVqC76i7n0cXIxgpnsF1ZAMtjbvWjgnmeGW1ts7mAPvtip
jWxkUuNtNJ5oAqYAfknhkLpC30qPO5OIBIIm2E4M7aH5n547cUyFWhTmASkrOeSQA06G0trGdO7L
2qCU5Rq9OR4Gj0tmZ828mVUeirDkGwkkT/eee22xxAS+lC2Vi39Q3/6PPjtrFaKX2vsfX+XQzk9R
Q9Nm3gpFeU71eoncRyhBeNPgLFynEyClKnDqlCP+x2cim3ItH5l7NAYi+8+Gnx4fJ3emojZmK5ws
+U0bTZZJWLWnZuK4W+BEeFRVt4IjV+XbmGMXDy+0QH1oNUKIH00LomL6YWD1hUH3U1YM/CNzpkS5
Wg1yVEjdZTcvvmgxFsnzSQ+XWEkWA6BccmBPFIPKu4F+yqCJ1X55ZlGmQ4MUgg2VoacDFCiQFKwJ
2Tu4IbQ/MSfSMMijyDFKRZeC74bU/QtjyLpA5k9ZZ0/9iSjEen+T3X3XTUGpTMys21RwZE+KuGfx
/NLK32ElGLFMRCsPKO4Y3HcFzdioErnBS+TrXF9SJnVvox28kFajs5gw9InWzuINSyXpf5eqlzUj
HR4MbDQQMbkh6r4SPkrjKo5K2DmOOm/xdsG0R1VYq/2fdv1FjxIOGYkUih7olDQj7XiStp73chyD
sCKoXbAiGz44E2ZQFkXda6kHz4cqdDN4FZbZHXWsoe1ZXwbR8GFg4Y9fsm0Aw2hVbocN+QYgHn79
cQ+X9TtpuXZ8Tn073X8QC5Dzn55z3faj6fF7uIFLUEVOkl4IiPcgUN3apejcF2+GR0VUGlY9Q3Jz
ZJJghcldeIYJ33W0wf15ngIyS0CKhBPueRcShS/+2m/p7RtyVoBN5tlGTV25/F5BJxSuCjndx4Q8
TU7p7WDbIipqJ5hPtA2u6vxf5zZBTG1lYfgJnPCbzMMfiEo42WWdgYolj2GFrJ3brLlmgYnLLjGJ
fAhV2dfOeQfU2QJqgXnRj3zVWr8J73Js1m4FDACk3IlraF9+GUwoGkKf90nFSauF8KhAzpcJtXjZ
NxmI/QIOh7LyaqZP9nnEbezE0DE0FiMDA+wX1nYo4wlbYS7CESGtpjTHu6DXcU5NfK4qcpFMfqIn
OJlcVNIudkqKf7rmm47Dup6hKaHHW1jY2fS2FEilezK5LpFDBkDgfsocY3UFxwICCeWs2vmOc0Pw
oOOHhmBbuW6kRRQp2ZIDD6FSrcre0sZc0Bc3W6vAFcYbMS1FmV/5eAwx+ZWiOQS031YSLxoVSLLC
6i1uQfw3x33xXoMU1Cy0kUdmgeASc8taQQ6TjSb3CqwtEXxc/YHnBpAyr7MBGziJggbCCJ5u8su8
6cZgG1iwXVXP0qSzQ38M1vDxhoxWlb0ykVwQxBKP4oYSuGDKP0JGFlRLfLKFwDXiFThkLMRRG1QM
ezVse7oG1XZUSqUBBO97nbdDlA4Lg6DRmGdRDUsuHvOraefiSvyH+rYouvCNNsJ+swF5LIQcWdUq
B7uo2w3DsCBKhDYnUho/7VPjRq9avSCTSZpcee2O8sCY/R45R1pAJWQj67diuvKt0T2WCrAR8pHl
qhNPahpYYh1NXjPh4rCXtkLp9LO1UHVBArg4iXAvl2lhUrGjFJE24tchxj4YT0KoVMDE7vEyOBGo
sx3W8unziGiP0WfQRCkExEMJpwr2dfoTBKWdHvwtGCd/QTblrMRXWZbq8N9bHJtZX55ZAjM/zigc
VQmDaC6GJjNR28OOSYGqTL9LWEiLY04GzXD8Qw6CLOfPRBdsGkEQ2LLqLMBsdL6GKazZHcsNhN+S
fo87vxdbP+ZIQPM1zWV0CN50O6Jj7IHx2xj3zI7gkvQcpfntf3jZ6DUhCtmr59pbok8Xlo5bYX/d
iyNdYySjnioKMW7ugXf7dLLyl32dvIUD6y9N5i5WXOcpOIJsbl1zoLAzKSE1a5m8xFd19c0DLUGY
J89ausEuIt5FVU9OpsoJDc+T5FBlts+gb17DqEWpPdrClXFmw+j9iqnT7KWn6fn9UQqXAoFarE3D
p+TUmFhNeDXrk+6aNLoAwAz6kPCyd04dZJiK3N8sXV0yDd2HcqQ6hKI1M8W6Ic0dUrTM6LTwxMCf
xrXC+hKHpydGiCtTHS6V6FkVjwukl7b+JixUnOwprHn/CAZNLiAihOp03Hd1EWZthLwTxWKmmjU/
bndKKPHfi/lwQznS7tkQpxJkTYNAQHA87ME8DhufYkn7bBhb9bsXJtyMgN6ufEl5WR+Jw6pHk8AA
IlulgbEeN84hQ8/h8jJeTBz9onk44wzaTG5MtTEdl147pWJ/1pqta5Pv8vdfylC3xIdwg0TR8c8J
Y8Ba0ESS0JHxJcFfMKqxSWStdGdnkFulBUkiYQax6v8R0zQfqm+yM8KZdWL8lrs3Pyf1nd9/L+Mr
aCEVsIrMK+ZMxIOXhi8Cq+Qhdq7lK3XaPlveDfHanD4F6mJ3SZ2FRsmSVvlR9APIDKUYLaO+2bkE
fdRyM4omfLtXpSffAmUoZLTsg3RYIwGKfHOyv6joZ6/scIbytVNWb0BODiORZ6j6qJ5h02h5lDIx
YpHxNM87I2TQrTerbOifHf1tvBgKG6DwcUzCvVez/EIZqy+JMDMzR4evUMzbmm/8Rhtk5dGBVNJE
HjDTQop/se+SoM9haWwmrLaMPNdJfcP1jGy1YMpCCcP5QyXgK4HkdqhYrZVTls8x4XVchHzC23pa
ft7YLaqQ1L1O9gG4Hp9blp5DzcqyTjLW7uSJdH3yd+SQ7oYHcDSE9HXyJDyBZw4e4ZQzXdvlsF5Z
RoHGxvr5KIuQLq6asP22o13UY2CqEjZhbP9CapspFuEmJWczctudjn1+pWTsi6YD9SRI3xjWnl8s
4vgzz1q65RQND3FRfECirHfpPPShgLnHfNfQuwCPy/2Sl3Xi5BQg78sfozAe2y2lpFxQiJoIgHys
RoZvimv6ac9RgANaJ8xGzH2VQXGJ47n2RI/u3Ek5Nf+PwRYeT0fq1+Kxk1Efgq8MrSLqxBW9lZba
Gwo4vol0OH1wLCEL10mAMqPvCZ3ssrD9lpKS7RrkA+EvneldW6nfHrX/6de5v8ZqQ/ijhuezQ0as
JQs0tKQ5gTsgkFfsgUZOHVK9IH9HiiAZlh2RhTLhCXdR0jdmr5xHUgD47y9cH1hijBzjznSIwTee
FzoOPDRM7V3hwrKjvAHymCG2Xl6mLZ0Xdo16vuEh20CHj949+U/uhGW6K4WeruasRJVUzfqGpY3l
J08DbG6BSSIH++GKMUNeI4obCy4wU8kp6rxtE/1mkuGmwfLkiFqBzE5Sr31BUdZh+B7dh31yx+cw
Rl27OTdJrgewB869w4pBZmmivEtFBmv7Yoo+Vx/DK3YbOsfAnVZVgaIajg+30hJB6AnHdGBaDvXJ
6RN/vp6iQxyWrO32u2xCFIvNshw+yJ5fxdJx6Q/1TRPwwJvPw7QlgVxydXxKXGXJDGmnxySOph2a
Y8eXQi0evPf1je8ltdCy+ARL/7W+0uqogcwzzM59MnbC8MVlXCiBZ9cPv5FzTwwKIkwf3m/ruwry
HZOULZchW04Hr2mdEfHVfLeIp427EraMaizmPEi0Sq7Exw80XJRPtgT0RVzxVk2UwI8Uad4ut46Q
u1oVfEmkN9AvZ2SEtlJjnNpRte9F90fTkpCCaEWKiywR0IRTmVml3O1A+5m/QEAbKavc0TbFhrnn
+JttfkIeVjZLdzJ+pft4YBAL2Z6EKtkN2gQ4us/fjI2F86NOWUrSzylTXCLmMDPd/U7ILnhl2y27
rS6xLlhovRILOyYGjF5ehoakjuEL7StTJLAWQRvQCTLP4CtVKzFhTX7r00nf+SoiRKj1knOvRSSC
MBxKt9HWGKrAFfasaQJzR+mDeqLG2M/QLcwNXP1lRoyedt69L9LLO+f3vp+0GgeCFFznC5zFrdwl
OiJXfmSgehs0MnmJmAGaJ12+SHtawL3BrIx9vveill+luYRB17D01Q1ke9YdXJnCciGIaLVsxePu
+/jLHRGAwwTu5wPsXmloSD+qA+9uYmupL+rdHQCsS6I7butUDK49zu5TsGdNbgpAYX5OVS4rrBag
vfRyOwMy/3vFZoVl2McwFBlAsiANpa3RfxGCaOJPoqxg9SqtX3+NuoGq9Dy+jvBHT7wlShiWQfA/
zUPgyq1w5t5Ewbl7NucLREtAyhw5lqdoiBWb25QSP8wit9/sFDq5i8CzUdJH8Kz7R8GboEG1D9Lu
pKJOhpukZi+V9Pevk2ksoHvDUvpL46jrCSVJ7DHUSnDYyICZnfKeUsXaLgypCkxRgvqla3lLGDcb
alVZXSvcYRMfQh3gnttgAroLNc3nWcqkhbbjhgowLJPOC+whiRZUh0yGOm3hGzXuYwV8eN1rTTiF
y2PN8W5WCBJtabfoFOKKonO0fUhZ6UVKeE++EY1rrSX59Vtp35lBxwXY/xpY9r4JdA/zH6nG+H3g
6SupIg4G2EmxvD5DuHEs83hXoGyGxfxN+2A5kb9dejmNi1JINpmqlscp8YaoTkRPWlTCif3dF3vk
OZi9kUJv0YZ5fTBZr2/OTmmhuIzTjM4EZWjtZE/dXvlDB3sQ4AVJ56MBV5rb9wx3dbpaVGXrQZ+g
DgUD8fI0jz2vmIV42m3M1ysGwjNETBWiubpITpSpETlzTZfYr2ypU1N08KbKrCIQ84gzxRSR7WYU
UHMWSi2foMm35deb28IFI3+29zNo9G5GaqaNHQq6P+a0F6Ayjbg8lZOK4SASNfw43VYPC1AX0CJA
nTl9RABphaaDO1+gqBy8Yp31XAh+lLu6eVxspoqD4MfelJAcYYFrish2XlGXL6GEzYSkiQApfiVe
XJBdJNiW+QN2fC9lZfweg6QqQS5AMn1eXJ93pIa9ozmxK59qN3w5RdPGkWjdqfWzJkpNMcFPA5sr
3CoBZ1JZ9h6Yfx7KOlPZPyMqTidC18WozHjZQVtZvZXTa+JfcxFZ7jHk8HqHywpBEv+x/TzUm/zu
/3kbc4jFK5kuuU72TrINJr1WhdOpAA+zPHvvZWiFoANVxB42T6Do3FlYPDXrFLvtutvDQ9vWYpI2
3mpjXzrqcSmidIJMhREfkVxx0BORqwdcC2q51rOT2cf0K8dBt/wJlonFihPdcYuZQ65VXjAZzlhJ
QpcN8TyUFJj/sWoRXtpAWeySwiyh/rxE+AWhVAY9riz7/8B6Y9lHvTNKBVyUi8z28GVuY5EDZSio
4Et/ZpYwow+/trKIkZMRdtdiaHHGcDhgx/m7ylwO4eNpLhaHN+eVYBanaGcgVErlIfTimVsYM3iC
Er45cQNJxjYEJpppELaLUvsbnOtTz1Apzv8YeIRtY6qX+MgMlMpW1im7f+2dssfeddM/ANZ/LWrB
H5Tk1ORIiSXo62sTfiSKWGqth4wTL7ktXdkpx+yKq5Gm59w9JgGolHylrO+hz2McNb1OCiWF4a/s
nYLwoYHfIx09NFmQeczIiWvtiOXxcfuKmIs5IB3zY3xYtJj1CGEZZZsn51s9td5S4EYU/lvRqArO
TtclKNQ3dwcVYrkH6AbzfbsQMXbt5ZIZMzWNZqEHjRym8U9U86xqkRpzawiICUq97C8A1q46+FmM
CrwqLdcTCF2Z95m6VElFSp9SrJtFgzjhLZXD9InIDuLPxHF5e03gDqcKxDaE/2l4vPmkhngrshIU
1q7Ke+H9cS6y3q9/gikEiFUbiyjb/rjadLu0J2jQEfcoStMzvZkC22VvXT+d7HMSPvs9fmJnHAZS
q8uU2AR8UzFUxzavjMlT4KZhFMnEl3JC1GY9NA8QtjAkftTP0CeFuJLijARLMMuG5ZpEoQMlhx9C
qHZjj4gZff/hZvKfC7aPA24hwr7BhKSym1yFkmqIMC9roHnyXGpaoHGB7LGcM5RQrZ5Gt+XLMORX
bx6LXLMppWc+qCvFe9vWsw1YGq5FW0mLoGbhCnMbpYUMU8hb1oSP4w4aLE86RiLTCdbYS8czZz3r
kv7X4dvBDdJmnQZWJwC3tDqdZhkxlW4P9xaWNOwYpVzm35w5cpWPBvJV/0df/D4VVq1dOAsebldk
FzYY3HtalN37v+FDy3GEq/dLtNh9z5C7Vw/McSiLQfQon5PCSO4PD0voyLpILdDsCbyWY0nU04Hc
jd+FReTxljK9ZhARzPtB9QX1qlackDt5EFBaABzEhbR/LqVAmZjZuDqNvEOF+aR9ECnVvgBqXdbz
PGKU5nrun+YjnbB2VLV/19+7NGxDTFgWP0Dx3bi2UboJAlgeaXL89mRg1cplmBu6tELfeCkM9YD5
mn1YmX8vHz564jtfW+oGua8m0hvFiYTo/Cg3cVEaanyq9lmJZ/U/JFr7Jo++2ffNNyDPzssLkXtS
hDvHtz2r/tKwrRom6+bFH2kfZUuMHh9nqxLdXXVNSHhNFreDhJXZNRHKFp6RR+6etY8Ru9HAVhSs
R6nmFBNK8i6rKvfSoxgQ4QL5HahQ6QdBD4lmTknxix+pGV9YuqxbacIDh9NuFzkhRoBROlDEWU6u
daZQMjMDzN1X1+lFHj2/Ur7yB5OUr6glR7CJ1rxGYaMsM5VdgYnwkiewj7yzYmchTh1zM3z//k3M
sOT2mw2fDGaywrGVwuD+HvPAR0v2LfHKHEUwzSi57GRehGffRFwhTtpO6dkBZzMJUg2DuN+1Gs1H
MEeByDxaqcI9fCDRCu+jydNuYhEvbtS2M0qmIrKupmm6UravUMmDIyHDPiUHTrhHKA12ZNzVCoJD
pVQJtcR9qlMeUBtxQ7Fjf7dvbb+uYbR0rbhZSAMxOoWEnl2MH+WD5W1pLDLKSzGLYr5LCMpGnfdt
39Y7Nrt//qwiX6m8IniIf0F2ftwZpn4RwK6oVRJK41syAlh5AqLQRJ8mt8ibl57j65/2hP/GLsUO
l46S2WG7KJ+T8FQOsTps0OF9eo4vVY9bwKUWwBy8O0JRomnjmDBiCAiaprS/7tJhyc6iu0RSrZff
hR2dIQwHXHPW5/+n7prRF/MCXMUSC0opuOMk+xfEdAmyR5/CBjB3gt7SStz+ks1+l6K9bhN5MmqT
OtU3UdGlADkWKPKuJaUnaZUMCoDnS+5PBoq62RCeOpHxHhcB+NkuRwtPlEkvG5ya9OKXtm4qnsPo
nUJdHVlDYKb6tUg+G5HJBCin47iaHXIZRpKP4B3eEVeQSfCFRWKboOGlhv/t0nHwLojwfqvzCOqr
4CmlImm/A+SqZv8JW5QZNzJ+KF7dqHKtCHfE9D54cMWyWyyfAEk6mcrqSPIQ1NjUNRs8xdwQX7Oc
cinEGzVYfB+5hTMko7Ox/g5L1o4s/B69Atl3mZ6XF6wjviTlZMuQyhQnbVaCNFTXUK9aS/4iqXFh
yDx77DrQTUysAoPXHNK6uu8574SXG0IA0scJGDjCVg/pPaB/wCiZ6voEa9BDhk4zvTMDsSbC/r9W
h8OkPuqxnNaYslgclN1aZfgXFnUl9Ktj1jZcFPoDKv7FSQPYdCoEbiSAwTSViY4lCVeoww6/yv9I
QOWfQcWxqWjNqbX2nmMjAAaoBRkv9Ck6GODJ86PjYDtuFNQU6ER2l1E/h+pzqA9Ex4pYQ48xN+F7
f5JTKk6bdMOgoxrHXT6fAoS2cpmY+NJOE4kHeaS2UMbiLBM5lB02IKJVQPxnGaxcXHa0o2PRn8Br
y/aW8kWt/mUuJ6W8gYGiElXuObgd4mjndwWaVRJkebVta9lS9GY0Uht59G9jopslwG0kFSAF58gU
ESLfJJ57g4eA/qDrC23tpJ0NCJ4IHUhfQu4wQUHb6vKLqdpH6/Eg1nZAQc1l25KRhSRNkbp+iNLp
79fOO+/MI8fmFY59/FrgbOTHa3NAJTNz0F7O7ZsNEnDzn58Dt4tBk6FFns43ZvwbDfNZED6b+GGS
QCQLsuv7H7dAGnYsxrlAoG+vtbWZdFqFm2qtXC3Z8p6rfZq+7WmertM+0QIbPq2JVlBqgrPxNzR9
6RJtNS3t2GFibe0RX+aU5KveiooHS7wGHCQ1sGz7y/Wqoj6ogp07tKev/QIX+iaJh8iKvGn4IqpW
9uOqN9gk7OBHXJO09PW9wkmcp7JTtGIBLCCTf6fJqbbbcZzmFxMBTf3u2bk7i25VO5+FnGueMfeV
O/54EcQ7Vqx8hRqWpZTet2GYynt3wNKEEWrMb8BrQaeCLcI42YNU3qn1GVgaWf6NEFkQQmUQ1ac8
v1QZ7eTzYxsGPKyAOwv6RsCLiaS6irt1g+cyU5gV+SvXfDPYDv/fQd7vtXn7QUuF7h4g1SeR6N28
YbODtsDbaA0a0AdZ+1mJ1A70oAYyZ2bq9oXeovk5LQKZIT00AiVVzaehc7DMfiNb0XSxePCokg9r
v1E7oJ8oYmnNlvD9AM4PH0k3ER5ESeM4A65ORPytmrJVWrwsFXB90GetwUM9c3VaeVzXJpYwlUpH
KyBznbojOMadRWbdomgHd2iHAGr8GYOBghrJM+qSDr9T4JZobBd7Kab4J4bq6NPzvDedxQudfckm
DiDHVGFEMyw1Cm2TtstSgZFL3b0X2ZG3hgGWTWhxHv0k2cqzi7XfJm+pm/pEu0y9DdjOFhJiPGIT
atFlDg8Nrmnjwj3PxKieVi+rIreinIqwgF9fieohTJC/JfHUnGhRopZn4oqfRnr2nyUpOQoXrh1t
wrnM7d1puG0a+8KKY5PEEKtsBcr3sD35nxSPwJyZ4DmFg8aqUQ+hfccuSkpFr5Uk930gkbywp2wn
q5cQA+LJiNwjvUrxPEfSRkqPgRuGMN6sfVh1KN7i9n3zAgVzqVDp/Ei1jAShVxlOiohf9zx7nTsb
1vdvhbvx4NQB81xqXqcKKoQyvRqElNJj4axnPQJW8XQH3e5uuFaAeV/B6I9lpKVhbzhIAL/Xaug5
1St9JX7BXYARMLsf6DnutcJFG1Uqw6RPjnBqX7OQVifXBy66mMiwJQ9Xoa6V0kHq6gEkKJ/Ps6ER
0N37q3EjW/DY7W/ntZXKcs8dBXLdrbQbaQlovfdPK5HT5a3ghUFigi1Sqydhk/yLwEzYiRBCEJtS
9JrMPAz1lkz5K2/ycv+8+fWWwkZuQONUw35rgeN1yZ8T6aYTi+A0WhS1+2X3oi3lz0p3REhw2/4s
mvbB+cLIoaV+mD/GOkzvmTeVoJCOp59pDSyw8Ymthv14Byx9SXvnhq6hzx/+BP3qCX3hvO9NKmO6
BVgerlNIXdpich2giu7kSqhxIvZtvSZpL7z0S+JbDc4yhxl+aTqczqjgvfMqBZbYg5D+rqbq6obS
Q43ch5lNiPXk1wQVFfc3PqwHCXde42xhu4a4zCrIiSS788G6y3m66Lrml2qCo+sK2FDWU6u+hBB7
Mrhlo8VVDEyPN5WmQT/TvjYRBXG7hSBodhSTiXbsaHI6xVaIPiOUYeW3Fvzo6h2TXDj8woSQgHll
6dsp6NLl09KKpml0h8rYDcOP2fOaXIIwkl6EEuOrm11qrBmoDmECOnPj2RWxfajjjnNJswY7NbDp
o3AdiRyXR26uw1j/k5h+v6toPOx8h0HKb5NBNlps4q+hvHKk1IP4nAO9PEElO8n060TFLw/98S0T
HZE78Bmz33KLLFgsP2IuBUyMfa241zo5a15T1U+m3kA3pW/3br7WXKo53DV6gikN6GloQ13ECivF
PQrMEhONttx5Pp+PEhu9YTyZCHBfq9jQhP4n9oc2XmCRhrtlLhKKnknlEugB8WtzlegG+wyKtiej
rY1dV+tK7+ce4oufihWHcNJnnBbMLS818iZQU31zxiYESX0sKiiJmeXQKy2xDO442XXmVEcoWsye
0f2tt6qe7Eaf1waignWt0WrcUQvwJd9AaNWJe2xROVP3eMcpVksiUKTON6IWGJ9IQgU7bGgt4ser
SUeGr+xl8GxwdbDlEY0sQekH5RKY4mBblnKexMRgpdDVgG9TJctOTbxY8K1lOTv2OxpVxtW1pWzn
kkXyvQfKssIq3exOl8BmOOCntYKNafuWLOtDU1BcM9V+rZTzUqVHdobtk/kiho/NaopVhXXj4/Be
me5JRJCro2D4sJrI1yzNm+8rDSPJYNouc6OTjJjEGiAJpiGdtw0gD4KwhkwNfhL9lMVHxf5oQv0p
5d3m/Fx4Fi6b08bDoxSOAn19WHDEJfvaSQRZtppOSVCYpo1pr5YdiRjjc0/BZp5WPpED3LQL1Jzo
7I9CBZ27isg66140xeeQvdKc9Oi2OOnPCzcEE7pczdKWqY6TNHSrXXWPhEI2dTuvq19RZpIQCE9V
7fAqetJ7/FoxWlnMQ4jrsQ8jF9jdvN7/TtWd4qWco0LEna4sWEAEqDA6WLdvU+IKcZKb4/UZVua3
1vgBTrKBciAsFXugCoMJrUGW58RDP1bSh0AihqhDHPTFIUc8An4IxpEEArD+ww4EPR9gbw8M/ZLZ
XmKpx+1UaRmi4YCAqaeyrZLO46kQaq4mZHuGXSpzU1jyeTM5L2OeHcU7ltocci1USVOnYtI2nPeK
zRYhD4X4KiL9ELIGIhu7LpWwfURlXL3QUEozXE9GCUpMn6nz2hiRrWBKJnIjyPNtOV5PSpfV9ean
MA4DvT27lRKgd53VX72pf+zHfFeByaW5Aq5VocC2RFYfvsvhB597/aCO9wcRi40Fga34z37Fv7xG
w/VU46njI9hzQqQYgs66CVffJYaEGTPN0T5miRKfEB+wc+eXwfuOl8JvxKZy9b62MZgqWCA2PLqi
EVI/bpNLi2PTgxldpN1oD0evnSwXyx9jz/RXFuiXFw5ECUjuN+DQIOg/oZwGn1sbU8fhkGUJPE4j
WFyG4cRS5o9ojuR0u0uYPpAE/QaD4Sa8z5jptBQHMeFK44QOGCHvmevGxFcR10IrVGp4Lx3Vg6kX
0Mxa7EsO7RgUtM1l7zZxMJCitSHciuQbDlJlJTAGhVo8JR8Aikbdd1WP8ObNljGtdvirgSNMvWsA
Ar4tRuS1YGH9GfCp+6Buq2cyhvBkAMVqOcNOL9ftfQjiVZngaYlB4ps7hSMXupqBrrTbrYiJv9Lu
nXkiA+bWfAsI8uNHw2zPlUCMr5Q3KgkLAraWUbm7gZCpc0YZ/wsBEbkVEHn+GyWCLVw40AWO5WGo
WrQL5u7TUVEeYMKkroMo/71TDiAr7UcPk1enLibHY+Tk4+N8zrEZN0GZhY6FrjMDHKSF5hHfhENY
9V2Hv8kdl/eFYeUZ3g3GWxxelAtJMZ4msviLxkJrVqQUxutpcSn4U2tlKY5w6siW75GNj54NuJIi
4F9Bw9yjQfIzwrexCPUQ4BU23viyksN49+g+7p1FSEMFCfWrxVEVN6RdDDRRW4krqJYNMOhkTW5D
Dgw3W8NuG+hGjgxGzksK17YrvVIG5tGDTJZdyF9ZDyVUJXv7Jf+O53tygDRYb4N8RtM7QxL3eSbb
XSPh9U+kcVJKAzcE3N6XDfnQzuf/n1vl0sDP/ziqRstkuAV/i99oeSgd5iZx+9LOUqotOVeoNHg9
XD8wCCrQ9hvSrABcu1t0B3p5tH/ruJzmJijweA4P8tcZ5QelV+e1Lc+BQORo7qozpydCzeMCyMZp
/ArKSNaJiEylEX621pLrQp5Uf6ROKvBuh5bWy95eXgaLgLmrnJtO7tSuYOv+2CNXbsksS5qit9XA
2ybemdkOTNqM26D3u3y8tRvPuEh4g5H6XkhlRp4a506/YN7TFoOrXFbHS1kbf5Iz1rCL5SN8WNj1
8kNZ3JfIR0a67Vlut5jhK7xu8B9RxjkBWr+ZLQTOn7r3WYUGdrLoY01v+mR+fZjFiKreKkgtrxcU
9kRIZenZPvdoAwEYwb/m9ZkmaBVJP56iLGwaoDK7F/LMuwf3cpH1BNBoJGmNf/1ZMQYfJrGgXT64
m51PwAFAoJbO5IyVmrQTrtM2xHO9CrDauQ4PkH1G88VMkzC2wDPELylMmGH+Z2zW8ahbzKmfB51s
ga17+O15saJ7wxOqqJLe4/rav7Lsn8Wg5q9L2CkEex5BDToqowRetmZK72KfWqSp055lmCINQx+m
ogzT0vkB6QBc7BqUWPSCTexl2A2KjNEqwlQnxAPJ3qB0mzMb2sZXHBsFuUPGg1HyhMoJMYspLud0
/Yxkbs1BszD58pcKVE4U/BuYybgKNndUMiPkNWmH5ea+P6Nhqk7HyUdT81vlZNkf5dhH/naQ0IID
NemfWPlEFzOqTF6dGHjhptf08UhISLI0UIypho8uirLDuyXyxiSnUEr4gVMk+ONXEmxE928v7YmP
2Sb84CB6RZeGMX2XOiZJI9MwSPAk4hI4YZZduKq35uaZqS+bJo9UkPjN+xcpHpdxfFjJc42QfgPF
vY+GNqcR3/SmQnE/9csBV7IkR4pZcJmKWz/H30tbgFQ1KghmdcX1KL5eRSyspR6HNSZwEqjCmDm2
cEF1OSsaE1PLhox2LTjut8sI+o+qBOX5HaoN/YOct8W4yNt95EX66VoUpIvdnZfxwcLexqhRcVJd
4wf3Pw8dpn0PvdCIfM6djnwwT9W3tKCkdVgNFmakSqGPPQY6FQ7jWXu1VpG2Rx0QbNR+OIAOsWTF
PCmZXIwRAVuq6tZ95NRZ6bcYwD7EpkY4NPwnAsiyySSa5vzsFq/LXHKMvEpZD9EEAktHj8+O97ZD
pUnL8pA4IGAKpPNU1aNfEwrGJup7pN+B/tfgv2VywoWNFsoGHET80VeJbKT+U39O9It6l77IJdnX
mQQMzaSlBCHv3g8yv/b0U9uLWGTBiQhvXWrCf873DV3IKUO2c+IrdahZCwTIjHltXIPode4xPhVF
TL6m2I5WuMT2ujgME0/Zg4yFm8qLy8I4zuybG94sBUOXczEtnR/mExsWpaZMYko8X2ZxT42Gz1PF
t9346sxA86CNZIqVwJjqiNHbLP9jSEtfKxFEyJ0pUC+N9tHDr/FIDFH311Li4tdT0cAX5p5irgYy
Xs31UQ4wjzAFlEiByWG0og/kEx9ZNrnGI5MuC+E5Q0ndKn4tjmmOubXmFEorItb0VCcdPi44UPix
lozKW4AQR4iuSEKsNy82kt41JjGNzsFXDgokBXXWY2m0X4Ek7d3//NFTBWL6ntZoFdSepQk/YJtv
C4Lb3898vCiayT+w/TKfSmbdboZbqqW7f0jeKpjPzucmWBgYpy+LS8rwvg3ttfvGErQePl95aUMR
nMt0vMNLcsEk8O5aXxmjkhyWmDukQ0Scd3ldvyBOVGEtFnVUmOAdBvhayg76EXijETiRuromtMIO
vjEzrnk3jvf3BKuDmUVa5xaKIijtMGC5g3yPpS7mgsPndUmCr3k9IB+m8ycVxt0N36XGFS52v75x
7eTTuJHIUudDnldUfEDnQbIs5ke7TY0MZfgvcVVCECbyhpiwUhKFtYkYUyMbNHFM0/8JB9EO0+fp
ofA7VyUbZZGq45qBHdAvpeXXaiIbshK0lbHRZEMS/CcZwz6Hhyc6Y9FK0RJNGNmQIlMwBGfwyj2Z
dIf18YmpxiQrdn4/ECMWyznMzPprvppxXUCy1ZsT2ryEjzT8Fv0yfP/QUFXFQq3IWFHhgNgTQWou
Dj21ujhTiEW/Etz2/BQPeFnaMikcjMLF1ytDW5RQ0ZL+2syIbseOX0oGrivcpeD9pvBUg1ULr1Dn
sraJHkSzYxkQMD5Q9lKKo9eSA97zVDU77WA+q3xJkset3D4eCzMh3ke3vnP0pNbHDQvqy2AD/+MA
AMmOq5pXvv2iLBu81GYkPGAj4FeBwXmCcDjFQNLr5myvw2TcRB1d8OoBkvS+qio2sezYo6PdtCjf
9jztXSlNvi3yPZgpJFSh3sFZtPUGmT5PlHhM+EKtK2EsX9SyU9Cv5U5a8tfY4WxuybIxE4LYMMa7
gHn5VZg3+9PvqtYLaSIXio9coI8O8zY9YMvS0jBOvcWj/Mfn+56kJPcl4+T7cRNJCbuZ/LXufSlw
wh82hZnFuwJssTkZARlr3+1VEa76X5lArIy/8MQeDBRFgb6EWZC5lvvpOtSvpGUQaIlWLogZdcox
Vg5KBjfJLbngOSTNYktdSOz963qUrgCHuQN0QhJ/1wuys68IARFrCtyP9mhXex29uidNGkUWqnML
QHUE8DnS0l8xQ7v9HtYYVlWazkmV8gQsi0HRtjbYe6l0a2TMhCJF1heLAN+8T47W1UPqqaY8GTtn
EnarIxpu1i8SHTcq+OtmQmTN8C7snZjECybqHudKbXj5XyVzCI+cvwvWmM3AwzmI/2vIrY6WWi7o
57vv3N8TtHFnsq6LvmGM75tiNHQ/8LE1LC9ReEj4mPtcENxlPhAA3qvpJPe4nXiY6tgz/HvlLUCv
Vw3n5tv+1ogtIeUUrgZ9R8MnjMQ9GwKPCG6bvIS3AIAWUCTTnjIEGxZgGT9wxpIYZzT57lJazi6q
mpK440GZRuF5RgDNPxD8CTP01y9m3m8SF0XRw12sF7pUdettwtbM356GlwrYWw41r30MRm07eKhr
0sXr47hzxCVy4gLqVQkk6lOZGpgqOTTTnuKkWVfpKu17dxkVmO/B0FJ94St3JRxnc2YoGd/5vZ6K
unWY6cl212uRSIwMo6O4RCbByQIkG2C8DjGPBo1sEseRzLBjpW4/WPiHyleXqyy4Tk7DMFRH09Cr
xTuP1al/Ifb70by2CO0gjGJswkNB0df5WTqpMK48t5vA+C692sEcSu7B8J8V+R6JjJxa9lLLIyyD
AGlAvFOY5C8zdWRmgQiIidWxVeAL1CuqDk3vL4P5bNo8oTW19O33uzwjN9yVUmgHjE4snfwNRXuB
pxCoc/D91xxveDJmLCH2ioL2dQtBCcLNqtBTsXVovOP9pijTXtVG31B3IhhZCWL2+bhSV8fdT7BW
62Y2C/4cXjB6jwGtqRw8M8awRlfVpGGMFwy/R94J06lDpzmadWjcIlIAwm7nvtDBd+HLCSL3TvcB
ZPc6waHtfoHe9owr8AN+813GEXPcmgreJGgkdOXS+JTn0T0GAnRKQEpclvwdMrrF4EBU3M3eAdZ7
x6ie8eqHQNpHaP2QRQYW26r30SRGEyC/12iKz4FtX9RDU3Z4EobFu5M2sR3duJ2NlE6Bh1a60Sw0
eOu8i/uuhifCzIBlIO/Yn+l4FuZ1/MvLMjgJBkSagQ1bTXxkZCSW0Qyg65+XdxP7UliOYKOR9Oyj
UEKv5f2PZyz+3xrFB0KX7pWAAuEjmqMZ4qSRQfaYiEqnE8VChcl8h1sCd89+ulRziZsUagDHy7MV
LFFGf5S2vvKVDZkwOymv8lUVn69iw5jPxxVelU/pr1IgOtWOUansVQUmJqoJ4C0nFJ7H2tUHL2X0
cC/hBglSeeyJWHO/kalL4KghfsHRGOqXefZhN2zePpQNcGm9FaeDXl8HDUWOVtCGfHNMfrs4uw/A
WR0g/wRzhe8Ou9MVSfoCJOzQMo9OiDTIur1mzPZbMpX+JPMiQ++DlcBTHMolBxgJcyZ/Msdhigco
TCL/mvgigJSezhz7SEqO8YC9EX64vc6H3CSbLC//riPGbk2UQU5EnnqISC7uX5Q5b3/Izu7d7Mod
+54gfGcz3YAjYX7BQD1KvRUbW+mwp9w1b3sVitR2EB6mKEmNYQTuZdAj1C4aB/CC2ux3efrez1K9
yEL9qGWTikQQ3UlnYI396BwzUH8CvytflsWuzvHMDOT3F+abUkpp/njpvOt9g37rXJmCdIEH7E0Y
iSsXtx2HaVSkqqyRSqGHXUbwC8pgkI1nCy2k5N5vYlUcFsqV3QjAMB7c7hg1n7MMQoRBf4otBEC2
UcqRJdK5qFwvWg9leVT7MdTMG4Ne3UBWRfhWScy26RPXzmNoZsK+CNG2jujGKeSUyasSzopknUZS
WTZy6hcP+CtLE0EUDa/I2L7hewav76OYsU2JH2M3LbNbhlkqaSzWprfPiOHMVMnoPo8wTPmn6s2D
xMpmkjHho3peoUWYq7O8x5xvmk4k6gJs3hYnD3k4YD+eseh2D/A0sWzNvwiKFsNvK+noH7IBXZbY
IVkT6cNJXnrrFwFk1POqdC1F61vfIlSLn+qVpwSEhdmktgQmClrBd1PO5LP3MpSNxl/ZpiR1SdlH
4xwNGHzgajgKZmiXdl1MLPDIEh8I1zAhNvj5A/opXJd1GkOuahmWfGChbdnR23rp5enT0bdBBPAM
fF4mCgfgSUHCg9BBCKdyEjok/RfJCaeoR+IMaYDa+m66784DvlU0/sK1M5DFr7Gx4hkQEScuZ7Og
5Qh0p2xxHHGsJoylokepzxvY9bDqL952EgpxjS+3XKxpvlcHtRViMYw5jKyaaGidnAltbMccA/Wr
3lrtQrUY0E3yy698gmNAnTFxNUjRhzwxnKVJlHDxBDFXXXKD4zIKze7Ln8oghGO4SX2Ta6yJhpGB
keFiqbdQXqDZ7mdReEek9x+i1saHdKcJuNR/ov7fcPC7pWUIMDRceBhuMte6UyBqVw6qY1Pm1oOX
2KCIJUq/6db321xtFmhwPFVI3y3zrZjbHH5KYcHXCT3oXqnFvrEbf3nSe0AABmPcLhsN5zMSSoIf
VNKFXD+PE8mlhfpBtTdGIFE3DoZ2abBfbprMe1J78eUS8oCIWNidyFQMxye7PlnfNneM780vnUSH
zG1TBoYCzGu+sLMZ2nU7Qc787Q49VenmJBJCizxqhyIBAvGYtQKwpXzxjgY1jIxB69KhpGcROJXv
sdxFmLkNUrZ7P0E5+G4TlYvk+P0iIsTX4z2gIl/ztWU8Ii1PfX9MsmKcvfRHSvjTPxVikK0zrO78
zfbhSKhB3XQbTufiwBX4y1VAgo/V8hNvnE861BdF515RjFlK27eemP/3Qka+K9z1m2lvA+XHytMm
234oxc/pBp3xIi819QD95q6DC0w401/B4dOnkk8MrVtVmajH+hAqXGPtxaWvnTKOUjDyfvNOksmb
mHZo+WUnuByPnMkIT+YOs7UsYyHFYnSwq6tyH+2CBJq1ezEpGYhoyc/STxAttFrwen4ueMrEVnUc
uHJXhnPAfeLHvAMCbhtTtgamBz1MOPCtawh+ZGJ9VtgF5OgxEU3k8nE3CLbVaC+nIf+eSfcfaayk
0ZxXSjBo4/28BWnejYxqXTZm+XkrNsppn+60dD5Sd/r++mSv/9v43UILUgd46ET8Q0LqGfZrpZYf
y36nMhhNeIW/7kZOps7exKYf72mvO2j3t+RpUwf3lNulHieDH2KgpAVnbjkQ2cgRLxNKnLpDo56C
mTlLzOv7EgfUHXfV00nNpDFTHCteUdwNh4RLauPQ9zUzPJ2zItyoLk4uGisLfWXvq6veNxgxFHaS
E1WAeB9NiZdEzhteNY5jMp3k2SX/wnp3m86zYSdnEx/ghbq8Wq3gBT2j9sjPYnh0IoJzOAuoRHyd
tqhyF4pjCW0n96OzJDB/rjUmo7ukJT4PWsWIMrDUNbim9et5Ka2gLz881q/RoU40225J5cJKoQQq
uXWCcCEE8gxeBtnImbuTzw4fSHmY77+iA3Ls6i99Y1PIfYPY12QuFSqPvLCgIHTivRRJTdYa0wsu
iXTWlNPwvSLMMqoSzTEiL3jiGSxg1p90S6sMj0oYjD089I/Wcl39GAqHnW/R3x3OIR719o0Nll6N
+pY2MrsXvSnHjZ0RxBz7Qh47TLjlRbvGmYLSQbInUlPzGfZ5uI7l6fCwh9HEDjouJELUPA6hVQIB
wiemO4FvwO+zvjxuE4CKT9GioAwC/nQ41V76qYhgNb66G/givGD8iWq/Eopy9mB2AXKGwG+vI17/
GDgHfmA5ZLAg3LEyD3BY2tk01Fyyg7Xoz7wjkDhA7DexcZkOxOoS99XAhFdU4jXNVBd9RojwhM5u
6naWXgY1Xxsi37qjONHVhvc+4RY/dC0nz+Msy0TM8Dxrkh71RpOkRqRetFnKPf3Z/wjpHo/iDdpK
J3q5oFU69AW/WqXtPCSsJTT5LPDImd+oGVgy8Lh9W9jAxdiMiJPc7NOPLvkQMBoC4sWtx94wwAXr
z/LNqh7Q3faIcNyORwkGXiQ/0eH4sP8f/CXTTg9tEhVap8zcu8WQhOHyibQYztDoKXo/NuyRsvZf
cqehdVyQTg3BHsBAN1UAV2J60/nho3dBFo0PJl4lkGo+BVUv+UuAzhFVgk5I14Yui2groaIuDuiy
xGLMiJOqbQO4A6ZXkN0RM/tkoY4yUy1RCRytgjkxcQGI+1nTFQ9KLQmeDzXpnn6hH1dz9G+c/Vte
pzwd8Qh+cQWVEWD7E2QELk7+DUoonZ9rROV8hTjLu4IvpCU1JTvomrQR1KRpV/T3UrMxIPY+3F0v
kO3gkguX0zya98MTn5OC0Oc3ekUi5nEFA24zd8Ei1ofdf87nJyQ25a0OEUUXX7NsA/Z0e/++pMKK
KPDaY2KLDLG/lgt6EoI6SdbLjLjiGJm89sUG/eJHa7XhKfx9Fx5dVTcIJCkpVVxP55j3oTc0sm75
whvTOl6+6frKaI384Uu4VewInIIRfqdiHJK2zqw5p9+ft6udYaQ5tmif99F+8u+FaGIiJDXMoh5h
sOXLHE4MSyBm3D6g8llJ3m0lbmZ0YTu2MSNfs30VfjKXQ3Uc75hQFa7EZDVgCstMYFELu5X1Komi
CPmQ+TXLLLE4gytJVz2kwW9yaTH6S5Hv5xryNPRTi/0m+eKC112+TpG20v8QgLVg2KI0lgdBaHC2
JvQtOtu7FMqQ+heMp0jpXwLD7Uuf2+JiiqfMgX4JzaP7Q6IzbPjdNG4j9cJVxDsk5T+wj6anqKpZ
4zpJl+03xjmbuk0mxCKcfZuG7UBtXrdwwaLAfhvQ97uotaTyreOqGg3UzGNUuqbv9GweodTssmDn
huk+4dHh8PAkOO1aVXmzj4EYnqfqTcYmiP0mp8hLWFWtxw6l3LMais8QEznEeZHm2EII9IS40We+
ifIPbovjtTj8JuZUX9x6U+jK97Aa6MVSxB4+Ts/bRghj2VdBy/ZFlFZaZSgFKAEFYWSB8q/e8uyW
MF+IAyrQAcoPE9VVwUDlL71eHmBt84F/Z9zBndFt5HmCvkV4kceQb+/SLO7Dj0ZOD2HR2rUqdtqS
9Zyna1Yze6sET017cw9qNgFR8OI1HXDRjkTypKUxzz6TvOm9KWczoQJy+GzgXGjam67UfIHYQjcO
Y84Fcx1C9CMe1nE2ewzNpSp64LfLErTdvdZ+MBJIwIPSmMgFYVHQJBvOxpEquNi93+29Sz1PB6Tk
WehPJ3LEKBac/BIyugOdzqfUTeDDVJRHw7gC9SfUIh42Qr3kvK4XBh/r72cOxn0wQ/MxUURZi5da
iefqp06e1On1blfO717BSKwv8nCm6VT8jCk1xRILHx8QCjqzIOGXlsWI0B2RFQwfqRsflsfpN7VI
nvjR6cKEQN2lah5o0KLF7PePnKVUPigINRqLbqwtp2Ff/GxVVGSM98AQ48BjRhleipv2kK2x7Z1w
JjNEzvnL1ZiEpMzkRJhHLxIsgdGGPkyOAv/e1D7zelw0L2OwzZD1XEkce0aSwQH6AHf2013jOfYU
6Rt7pIu8iRp4jHQSHlwKfUv4E/eblqUrtY2T/oFFoFLkm1L/P+BjTC4jCxCrfN72hEaP2qNCMQV5
gKS54I3Xp+p9jwSNJnhV7KkUK5Wfd0EmmkpiEt+atsVLvtEIEIzmr0TKqR57fih2LsMjzUKPMujv
FcPXBNhg4JaAZtPsJ7G14ysluJ5cE8f+ONkpEZZXv3g5KsGed8EbcH/3D0JFkoBgjOzbai5iONk3
7bcgxZuKpo+LQeBYzIbCECqNsjqufdiMQvTLUjPWZE6E+1qjDUwBq12iDUHJKzQskXnFfzO8Lgdp
YxyksaffE+/3c9/ucoiVl9AsFQE1mATTkEr89aUJk9T2ncvrFMY68X2xf++LbM4fkmi55IwlldYd
CMgSEAuRQMoRGZpq1nr9zx8tt5le924o8nsZjzxaDIzpFHS/mvo0ma+iJo40pk+eYdAgLdOlEZzi
kB3UC2XCY46k8yYM25hXMioU/MDRJZYtQQ/L65uRVDrgylQYGB0Vaip+PXC3rA8y3ZQmgJP7AlWf
neKCtij4eEksM09cjApcOUUyl7hlWDs88FActJYZ3+6YEJPMrUm3zaPNlv9LvGbOQtcrx7Ii5uyU
AGzJQhAeyfHa4+3aqYmMtnJM1bi0/FBMly1EDSAx9o+ia5T2w+UfBqA+VB4oJ6tPu3xo3k4xIE8w
SUnnc6VTCepF02pF8CT39vCRF9VBlj8fxYSSFGseJSnfhRwDC2gnZvZpcrPbVfUh/hwhlmbgDnmv
9CV7e2R5oRS0q3WYurwM5/LxtIwvn+iqEBOeXWStX4wibkMWafqgqRtyZwU5nswHKZbqziSZFul/
EI/Eenuy8ngur/472LLipSOgnNwzRJJi4FcVSXCs7u/+wExbC8Yhou6w1ZDfs9Pff9Av87jVglEL
lIRuLQV0UfMYAp+pxefiz1jC48bCXDOB4Yd3U4XF/ru8tUpiG+V3E//V9a126BQvDkkQjPRCbdw1
74+RncVPHLKdXU7Gy56yQT2L5fQ3O2GRCsaNngAx8NCJr3r/QVuepuAcR2x8J+QkjYReY/ihDZVS
qlMQB5/WeiwQ51mvege/VAMHbM5wAbaAlywvMtzujqnfr9A2Sq/BfqV9rh4Gb4pEIQwVnZN4Rg1F
43daoev01OYmji8Z3LdlON/IO1PsjkEzv9HJMElPW8V8iuqM3ykXedz0d9pFMGYaGyuagRDpjwod
wAStrENC2O9yiVxJm5JT+PSXTfU4gJKp/rkjvXzK+D40j8HPjdO48Tn3/H4apCifAVsf7SltmEHW
bmzYpZT6/cUOlI2uzqY2WR2MgRdk78ysQOdAuDp0V2uDkISlroKT6EE2/K+uB4rD2CVJWFPG80lz
gAv6zaMIV+w8SowLsg1ihnAWhsrvWYJ3SwacGQr5TkatLRJnEBHRKeUqtcfFF6Pb5AjahLJEhjVz
j5yeJ5swOYurqPQO237iMr5aFmEohqK9Co4qHDxCNJEnue2F8/pCMYqLMRhPMOYVZ9qtAalVe8A1
5rVWOcKefauPAFLvw+w1Vdtr1EIIyNMhfCoj2+5il8UbnHOYnMLOpgKaxzPYAQ7IczMo+cDIdkiL
3aIoRvfI6vqM79es0PUijfMhpEYDc5hP0xvGIhM7e2VSw15Q8VLJ5b5YxKx36/D1rDzV0GDtIPIK
d37mKeVEzNcCI6+q+72zrCRcHFcQoMHLUy9ipKTvuf7ECpbSJO2VGm5ZiUMd+JLd5CVE5ceMOn3J
kmZRYxf1sBw7tqUkHOHyELSSq3cOzFIeAGewZUBGWByIr2os55lYsyhXRv8cCaEtm4K8WWUqwNvU
bSmwz7h9keovWIYEv1WMbV4FzYxi+KIX6yL+KGli18QdFVFwaeAPlh3TjHCleB/oiKSCN4HoYp55
HNVyUGShe3Bm4DnK2di6D3lJT+WfHMJwd0wWsDmLxMPEN23Q7IResCLb/kOGO9cYzxzY7eAwTCQ8
vL6VhyxpKeUZYIa32JDOkIf6KwMLA87W89vvNqPYoqf8fhpb+nlcZFzNtmeLbQQVl6Enab1NU+jo
//0Gocxy2kQhzJ+J8bljXLvkusDATkTxk2NYjqqNR2aBXFOCYSalOEkggQSnCnsNuYr32gsn8uO3
VLbZD/1qjc92jgIGYIskzpp2N+71F1a4IOwwFWBESn8DrSKFKoaW4kVzCzo9/MaXsdb6NrMDIzpz
hTUgsj1N0eIcJqa/Sd/OYf9Cjrgrww3NMZ2VJC6x5c5q2CNca9r7vZA2rZanuh7TMW01fYoqo/qN
ng/O1GTyj4OG1aT5wJPEpnjNRgaJHO1IUPh4cmh0bvRfNJ6h/1j/7JqWxqJQxk/xk5bKM6kBZrhO
uIN6K9GYvtbHdCQukr4y5UN0SADoIBZmM3DTpIRBCCGc5hngJqqw7SHz+8mopeWiCraVrN+1QgI9
xzYvcIfO2nmfTQcNQqsNbD9ew7XrNg4pqmzUv4lIRemFlFIVhCqAYmobDUJQ7UgzaIjvnpB9UnSS
BkIVMgHALKBzCXNJ0jBaPhJt9Q2snd7vezqlD3AK+venSr/f/uoVx55OhyUd4f0xeadsV2vWO+5l
pN2aRDRLbMy4XC5LHDTBMh1UoD5DcmwKX37/WLbFogmR9pXij2xYMwW5OJuLJw2SHYaO9EG+8bra
tSZplz26XC2+KyuGAssHYZl7gvm+VgvYcKMOnj9LQYAtfIg6BtU/f/BC5stwjIfmp0oHG0JuO8uX
3ACqmz6C1gSKvveUY/M7PND84dKxU2UHfuZ80bVEC5gKTUa027CgE7b+WTnmdu6XE5TSf+tbsH1n
HSeUqtQnHdXAn2T1bEo/ADVz9U9p/7Wb0VJRlDsHobTFfwPw8GcgD7EN+XNUe8qKqbNMFGMIcwb3
qWq8aA2g9f8iEtmYCJymQACCc9y4I4shBFeGOU1nDoaUhqk+8MK5bjICw0hpsBL+Tg9opRpaLocQ
XQApvFgnpNl8Rk12lpTOvQGFAP+H3rcKhtCoX1MHQMezqzW+SpdtvX20CHMxt5c/RO2HOI8PkBQb
WvWEBqulLjd+Y1ONAp3jJ25iZDXwOpxR2TDhsQocLXJoQ0shREZG3kFLh2IIOt+UEXfgRkgnS2qV
qxbV0ekXbkLzf3VjtjfbQmF9nPt4YSln3HHLa01fruaMVeY6RvMU7lNcn6HfGUYrgI/R7k/si0eW
0tRd1z1xre3StB2sYXqt6URAByo/krk7lAhcYE3Ue02ztmNNs4O3mVSbLPLAPTzqA4mv91/RaMGa
wftNsJ8=
`pragma protect end_protected

