`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ER9UJfRnXORgF6nX1AKUL4bEne/LZFndctkhWCPX6wqHo72wgQVwNm+P/rTmRg0gzsvhlVkiZ/eR
NGnRzuV3wq2ew4+ZOqxWQYi5NxC7S4aqA43ZhMdDiWH+PnEt7kXzTAMg44eVVJ+v2kodj7wZouwP
1H28tXD/Vy/sc8r6hpybu5FUXHFz/2RfiTcqEHI0RA5Bw5kyTAgrTTX5o/bfAEM2Hh10y25OyHJ3
vEaE1fWJDrtHXpYKkToxTTYKS0oInVvxqfDYHU1VQ286KGggKkj246YuceJktFgMsjzX9AdVvEns
x/WET1Zx6Wq6qoBEX5J5PQ0vig5DBBKjIrFRPQ==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
ZpHdnXfuAgsmFsZSnNzqRMWD0NELhulq3a/LUlDNpPDx/6kuS1GRJ4Q/oqAfEqA0C9hdiTirt9be
lhvJI2KW5JSVL1U3rj3t0OlQKxY4N/8/TxiC+e3DeB/QsXknjJnpoURVmYtL9xdLVEwaRfYCRBCi
MEsHrm6AJ13IGwJ7AhNeOF1VZq4La83V2jeZk9bByhyGz2u/ltav0iktMONvKTXtSHpHI7IggA2M
2FF7XLWRhurSxaQFQ+MoNF3Ts8wASu7By2sr7HG9QVbNYmvbicSy8l3YwKzBQ1i5ihkW18MVZR7U
SRwR32OMrjpWWIjSpHFEJIBbVnIZzpYVFeJMmgAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Zzs/OsHaxftOPQx4ZLNX+X6Jlhnis/mWZEQraXvNSCnGqCo3Op4xeIA8U1/sn6mXGOHpEgf7fQd3
DmJNU11edA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ipkd2bqhbdb4wYF5RzRCEriZLYoPZiScQ62AI8E3rFIb5iTiPi0V/4bHUjgA1JSvtgijXeePJn33
lFI8q4sHCyS/XOrgje7fA05IpaN1+uPedjycAjMd4AZFq1B32n/x+ksc0pSLcwROK0g23iqWIWWH
9rF2DDNIO2a4L4oi/ff9OtRstv+oa6l0n+WEZZkciFIWRX5EabGfO07mWd9ERCKsfPEs/ShnYeom
w28oKrROye8gkH2/uK8XbtrOuzWwBxTfNFh+WIpwrHFDomiKXLF/cFt+l4PU5swnAupTE+fRI+66
oj5r1CP4fFcpAlrdEiYjq8X3g8LoO0ybwBMUhw==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
h+V1ZN3Bbh88CAc0Ns3Boz18hwEn0WF/1hwMlbEh/V/i7cdC1hLjxC+5rqbsZ/AXnpvJxSAVwVwi
Dq2OPqzUCcik6pmEy+nP5Q/vM209c+ibleSGqA4dGVxQxtxWUtweTQNwmrYi9x1qmYm+wKjp3G4/
RWN+pvRQRqfkd0M94vjsHIYt4edry1DmBKVtlDBfV7CT6YTAK6N0wX8E4EE7SGZude9ZvhzfmPiT
hS1IXzxFwU19eWrQDMQDz8CuT+LEl8Ti12Gj/6iIC0ng5VWzpHQfdsjZUpdUDqu+IfOr2w9y2xjY
cqHmE5pRYE91BjAp1yiRiC7+5QoJR7WDM9/xug==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
D/1BEFzf3Dn6+qKPmrwoZj9syK5lSSYFq048R9JcfSuvPtCVMovgkfw5mM/mBqTwXoMe6ANT5gEm
6uYLLhG8ke5/TM9ysUTw6CNGZZC+SZrX92tMX+0P47a/hZhKthL7X4O0wwhOqy+PwyaybsCg0A3b
pQaGIaCmo8lUlBER1pU=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TpNEfwE88dpfngWeziW+u//YAUWQ1HXGxofatYh6j2xs30iQvwn+VAgYsINJqSOr4/VMsQGV4Bw3
IdaeL4zeb5rZt022Mzlw3AKQrlHGBMs9kCCytIyoc/X8A5+F1wUlEO8VZ38KJPBYOveixG7B5vxA
XrdIEKcL+XJn4B86ytkQzeSOoWFWNz44woaZ7YCYWRYNFMrVvIPHBUaKfsnL7DDYkpFT5suDU+Je
ngOkRge1/67q0CFG50xE/J6Q5sSom/f6BUFxRzZUMKtdBgDfGUcd3MxsJZyvZF12z2+t1kRvKiEK
OC0tw5Y8FcF7u0ju6CY5vpscAejXLjFRXVvX7Q==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qmimsPBs781pBccDrLYFd+JZdKzeZBAiAebjJio1m56BO8aq24X8vI8SeIFlq6fHQKFRKjlHOdXh
5m/KSLd1VUNt52WPIrjNgQEvRFcrtBuHmGD8rNpqZIOFKL5HiLgyJvLpJ7O+BxxSyCzs6+lx3Y3d
koRAF6/DTqVe6pJR0/ijoN3Gf5LmWWB/zfPF/FSpReDaTabkJBczftODiLQmSlVjlRl+3auS41aX
fxNwiE6EbmBw/AJvf4/uq3ZMiimIAR7beyu8I04vPZ0qXnmGWai7Duk6IhyIviyycVvBKdz/O6RK
we6ghGDnwxYByqw4Fo1n2u0zLPvSqhgk36FzJQ==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Msj942En5jfWg2Gjt6FyYAShYdKTfBivvo+K4Kw85jq72BwaLAgt0K5DLjW3ZYH09y1WrDYM6AD8
7gv2lnlH3m4gzZiUbWUnNPUWtnrDD8GvnwcyecdBjgWqdI0KWE5nRrnKYbNuUujafEtWYcOYr6FM
+26WMMg2gzy+E+Gj1TQ=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KwP3OO2V39NoVOMbQHtMwhD5GIXqQYRM2+ABg9k6+8a+KiaLQWvHZfldZ/lW0EmV16NsszJrmMLV
DUxXJygYunyrA9X3fYYcD83t++204wn0UhzAOy6QG0KzpoOf4oW79eOJuB2FZpTmnY9zj3KPDAgS
X5iEzu2gw0AaHbiEFQ43NlpyY6sObwn+Dxu4shA8tSVQoOmh+lukvVpshD5C1/wxyEOSnhKO4IWl
/4uXlY2E7i+1NTteA+fIuv6JmjhWEhMEmJ74C66UZ2ouq20t6ca7oxRJbhXR8+GWbgz2vHBzAC8r
FtOxcbpxoi+AU1xbQz2ZAFrwg0bm4/hY5HvY1Q==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16320)
`pragma protect data_block
9laBfExh/reBxdYS82RZrwLWqhPdX7czJf9DiuDus4apVEpg9+rZpvFsQ62RMKdYlw3hdiyNjEU1
J817Mcwi855bdOJ5n9Sb7BbekZUTFEsTVFSfC8xv3UkKo5NRb+Zjet793sBjgX9QNE2ObbaK0m7/
GOr+Ub8V7mbCYlsnHS5TI4ha0vpUKlyvcCAUrwSWv99FV0Ah822luJT8ifzKnDGcVfhvGg5SBmjr
HtvjEEdNsf67gjg5dcO3qVNKurWbIY257umdP8XBah9mCcR33C2D/yW2TFkBcWn50Ihrb6GB5kHJ
d+GN+VfyDM7Wx+yEbv4JD1qKuFez6Y340asdxCkT5OCw9kmGHS2Z/rzZzaEiZVFBy5UY5x3BZ3Ee
uXtq4tdYZIGdFQ3L9gJYfRh8Z/6AT7EWgn+Gcd6ZNMuaPq94ml+UFeDMvXolhCTYST0ZUu6dLUb4
aDjoRmUKfnRkWPxCxIXkvBz/uhx/ZbMkCrJEnbOQtTftLfTCaczUv4hahHsEclm2G1GSI4U6oOu4
nsmdaN0E8auUxm/M8ryqi73A5YrAZieKKCJwjOLtyaWz6nk20aDRa42MsS46EyOstr4vyAMgaVez
1njht7cNpFtaeqymJnvgULw9g2mYM0u5Cy1G5guJrQQFuVrHiJp9h8rdIuRAG6Pe6GjbRUDCr7vI
ndzFMA4SGlr2UqiZvxeI6L02Cysw0FZGPjtvkN3BEGWRqXuDodA54ZHRgkDLrg18HCgI20yYekI1
CtYnUj4mZHPO068TapPXrGQPbXhNSnfYjWLFzeZx077R5egEYx8BawI/Trqsli4qRj7zDmHg1T88
Wjmjo6VtTTWqRUM4dK/XtSGxpb9DulOG4WU1uc8ycBNygDFSNuzFVXr2Yea3QMqFq5gnMNf5TSoJ
DuNaMvMt38YGLuOS/MTgehS6Ne34754egvtJmxKN09ID6eo7RVzN0EpEqrLELfGkNqIk5DIh9Z/U
5cTJfnLhVrxYR8rK6PtvGbkwY1dSHNl3UY/p9xqVg5ZZDOIYAsUlKi2PNca9P2OGLKLapIJrCUa9
lmB3VZVrYnt5fs9dw1GNSKQQjp75lvlJCjtc0IvNGWjMiY1kDtnV9lcy2Nw/Uxe1VWj4Tz0MUfg6
fHZgGvXVdFX810R8ZtyGYN+9NQ7mV1cHZf9Ur8F6Ot1uLfnzBE5LYV4kLFJC0uYzOapExVZ3D3D9
WBHh5sfe3ewRvT7TG7PenUcrEchVB7pMQNI7KLfx+WDyJpJeULsgkbwQJZli8ANTz2Kcmz9qYLhr
GH2WntJULlAoGvqPeh+An2R16gYPsW8aiSnEHHWiK0GhKmEkHo+U1Y5blJFyDH5juIMcPPuCxtbw
fd8ulOVYh2l1vKbD4gFyww0UaeUv6kFU96JUa5VvW/hIf/igWa8TnPTacDVWNug2BUVsRrDkZ0jC
/d8c+XcTEMc3DEDnOwM8Y8HkW7ev6YdHejXJydGgmRXCUYYzkN/+4AHk/zhXfwj4kOUbc1Zf8dls
yGr5YgYWyD/jzcDN6yioU+w0PViTSDMY26VnvBms6/R7dS+vE0ZvcYmMhkr1dsSkDpVRRSw9TGVB
MEpsw4Tke6xtqTEobk5Odit8jsj9xlTh2EVfXZNTtSS19MiUDqttlfRdb2oj5zlDEh+YaWSIhDid
RVWb20bUrjcx/0pUlO2hsWWk+OS4oSBPXGNPN881XZmvBhOnEj9fdXGyo3+tDetDtzybZjQ6eEUm
rMmSp7hNPEPMSKuGjNNxe0xrXSgJ+EqHXA+eQ8N6d86y+AAv6fLrnjHOMws9bBnNtGcKN9DoAU7r
5F0KK5rlH3muswvXmNp0hjttrPjGmt91HTEltuzXAx1L8NqL+bBfaC695DdogbL9f8UaYA1A9zhn
dBJc0i8et0cs7lmzwk1Gd+icmmPaFl8SA3h1XFYv2uNdWQ526WruKHjkSDRx2d6zextNAWz8PPr5
B6z0aGz45eM0Rfkl06aamIwW/+g0wgS5Iv+ZFEItVRxzpPA1JOtF2uvwX7WlMSQcrXm0otM/eVQ0
Iwmrz9xbtAvaxDnW8b76iTL5dknSrwuQqi1v3AId9bjzEt9bSea8VevESn99T+YPp+NapX6GpF5o
VMkFYxWWUq3/4kiIw9inOZoSCQW0sWBx9nwhlWN/d8iRG/p6go62h0VX+/iC7c/KqSvt9//bw8wq
tATcfG2tZO2Y0SLf9UnIww25sJLNGwZ+MtNgtQElChgGZvONGYgQSfVuRCicWGQV8Pr/VNu07XwH
cWTgLlLysqQdxBbU88umhPOT0zbwNyyRFbCKv+L6hwWysWUWf8//LzAmki94fMjbmEnjBDKLi4jB
ePPYF9WpEU/J6GLJHwJHVWiKmxDKiJ+2IF/ZbFzp76EGnXISq3A09UoJCwvQW1/6jFip2Xuf7TXj
BhBgMJ8aTsCwDVl3dMnvXvcJIUFQ5utwcltgnAs2KIKDRhLtBLOuhB8eZhaHrcfI3E12SC/OBx9B
GDXKG9O9vfvgWNXcinL/j1aj0umadXuL4VLrQxUDF4OlY4QkDgfUBUW4nOplAEXhh5ZXdiNdPROp
QTw9kAIWnaESRUJg08ppiGYhu6xP1BJsYPYw1fo2XkA6dtIiN6/O2VLjWNIcZRrybFl5KdGkep88
iDU8nblWSr0j6SQ5z6gi4qlpiaN6IGlRXiS3aGvSyXSSg1i2lX++YqGAxdiqymw7TLHZlmjGwgla
jPTrETQYXzO7e9vj+mVsXvMjEXicDWQjcevUT922ji1oU/X+6RISf7PlDX2fwmrE0QbyEU++sNpz
l+gUPG5/Y+A6BnCS16HwBMs+eE3UwO8hmAvdzuDVPujLC47dXWlU6Cvkys4saYp9eVME0le2b4oX
bWD0W+o2si4zkaCVod4twipqVdccKW9QxM/V0JhoqkPnY2MJqo/r3uOKYMUzRXANUuoAjRhXQgBN
et7IfS8oQsdBScmDVfEQNOfGjzW3jFpKrzMgsL2u//iy4N0JGfSGx5YLCVSY4QT8roF1Hr0wurIj
kgb+XkEhZ0mBTeEAnppL0rN1opH8m0NNWdGrih8nUfpzd/ODSfm24WcGhlUGeI5sRMtiA5F2cknT
vOnHDurXQdJmXgiVCZTP0JuPqQyKdI5yE3ZjTxutWQiHfM7TsEdb0hztf+LBJj7V85dwPRiCVvaW
41CizEInTpeKt2xNgZyUJa2xxqZzV9fVW8pR3mKr9/7ZNKVjccU5zxCMHQUOc5Tnc5vTmxf19nMr
+L+4MsX6XpGZnmgU9ep5IpKzXTzDbfi8ghPpsZjIVpIiRqa54ga0xDaIu+Hjk/rLApFxiv6c7BgP
5tfMc+REzxTaX7eV3RYJOWtgpzk6PR6h3HkcCn7uIn1zhBDcPV/gQF1ze+qnCajRDor1zg5o08+a
00mugoc+VotNANH4xmPXDjq7vpaVKVu79aZ/45ZuIl6Iv1HX5cF/Ejv9uI+wbqhqOIGpPFYl1Hrd
XUVJH/vUT4yRV+JyFUb3qSh2W9D3fJTEgUsbYIB0swSHf3AZzKdKNZPsgdJQI1Dj5iuQWl/0kt9Q
KVvH/RE/IjpgR0w4dWEnO0UkJduSl54zyNTKdVE5D0V3bkpvQSxMy3FxjV8Xf5P1QnsXfa2JMemT
aw7Sa7mcLs/8rvn3yKyod0sTBVKbNsVSGbIYOYZwifJaGvQpLv7Z4VdcMqMouVsNG5kzT6a4u9V+
7CUf1JfQl0mvryDOrPrT2tKuaAsaQQTW46OzOtxKFCXtdsnkRATJhmzhUVFFaYK41jbhI+NFhIBi
u/U4SJdQWpv2TegaV5hS3IS1Lk99aTOdvbo0GquBjhs1P0ieBOnDMJe2ODubhMGMEFjxeoaFzdqw
J+VShdX7REcGhSn6EmiriE00kL+vq0b8UCLb7H+FAcF6PPVvWlgYdotQ9UT4PzmOZ7XfcViFzJ7V
ob0KOuO0ViSMEtVfISe//bpZ2g9QcLCU9hJoV634F9aZobD0TqCBfTjRrXKSbT0/SmUYPgWzznbG
AemLpGDMHHyk3RiDq4IDAFFiiQkfMhrM00u+Q8fagz8CC1uyqt0NDUbqt3REiEgXqHUir+VShbdr
G+5hB1KpWibfOoJIQMQ8NQ074mxz/kX7/K5t9bCdp+lzANUY537bZf8lymvQ0x/tYLHb1Jb1c6Qt
IQ8Gg978QSidFe07DnlMg5yuySA9YfPTUE3KbiHMRGzGS5r7qlXRWD8Pm8pTOq4BFW92nMxPPZzK
xqbWmvo9KyfNUvT9LgjIA9P+spYGPGgRSe6HDlFJ5WXYBo7na5vBgaQc/jeozsCAqe62qsmXa6cm
jiGVj6IBYPCfIk1ZxfbkvL5qmEGcB/CcVFuABTNIOMplIsifFYzo+cfIGR4cfRK++KCcmx9H/ySJ
JDvLfLGIpMw+fCDPUygel2jIdU5VCnz+cXtV0O6DqBko0sbD7g+AnldXvSey+HK7cGsqDlu/rBKA
b1MmFDg7MgzHDO7+cBAUouxSC+GX0SxAhM/35xMXX4iYOQa1u2doLFygw3u68+6i+2BmUkgabu0l
pTimkde0bsVoppFgWtz95BXycYyZ3ZpkImSayq5oz/fuWrLqR0deJ0uFC/gBuH5ZFOJrb1ervWiT
lSo7IAG0WKl0MN5j0pLTIenBKEryhRR5Dsx4sv0A3O3pJhLyHEeDbWyLWfgLp5Ru25s1tdY3VU8w
zDakP2U/b2Aa1e+G+++mniStl+C2ghQC+lxv8TObx2Zwvv68p1o+c5aVEMR1Xil4vmKfLLA3EHHZ
ai5PsLJlNd3qEHDCRgEUG4W6VIzBw6OzeB1SJU9hN584r5nLqDj23PZipwkI/uUJR9WyQWGR/MN4
OwyntIkGPgL1u4Q11x4zPUerqdNOgvicnjM110DGexD5XLqVAUgPuvUMWAshym9DjdFD80pVVXhK
tP0L44FPTjMdDNgHMFyt4AMG58oTqBJry76WcBLxCNtKieSfge997VvfPFoRoG2eq3wjXjT52H9V
ZVsnr0Xqg/KM+7TGkZ0HsMvKOL1i0/Afj+nuuw1cph7AiFQqFDx/3WbKhUgp8RB5CZikTodqJ/k/
7EtO2bIw9UmlBboMuSvJjWTA+0KEqxrCbQWHQDnB00WII8PGjDqBAnQ5pgh9v+ls3rp2fRof4+bI
AE5sImXDivWW2a4n/zjRMwgP5EbaATn8SiKRjBa/xVH8Axc+p5elUIvsX2Wz5Xsn3h3VPDI9IsK8
aDPRl82L8PsG2QNdZcKhUGxwOpTYia74HswplFap12sARlYzQ12PKA/t+txxZ87P6jd7hONatum5
MWikiUR+n+ZMfA5ovye/G1+FGzchNIUvEb/+y/Hz9pEousoMrRn/ddivdLAyzsgoDugfN3RYZgCx
lIO+m1wrmaUUgq6FpvUKAH4S4K7AC7Z/LknHXZntZGie3w0UOT+EfRFRawsdrqvFye6t7ZlQ5hRP
6GL6Us4+JzxczAYKegHzJZuFzpZbIH7voYo5QV7Q0nDz7aWBzXDRVYElKqtncDwSNO6wcZeU6P3q
kl24t3PqRTdSUlYLjSgJGQrROwWjC8EXXZwY5pySkDGl0BIpfIq9PWH6QT+hgLDPUxoEy5kHd29Y
Rsx2NvakLM9UX+TTzQNM7eHt3JV2EdlWRtpUuI4WHYpMxeakq7xoHSNsaiMAO6bRcthGnvX8k+Mu
c4ytpK95t+wDQYiWb9ghz1zqpGgZmLzEoQmhSfzeu0F3j9zDg0IS3AoYOphxH2OhjJoeHSPczSSZ
SYLZ6K2hVJpN+iIFJfHPVruACSImcSYLJAWEFKvZgCIHPlDiou6ZDtwfe/siQLZ1zZ4FBRA9ReFb
pODVXwlO49Pwh24Xz8xDHpRC0fPHd7O2ujYwLA2AcLj2/fCVzy4zvhBBXNvSAtDHz/vg4Ivv4qQM
xrkoVTDi/14sjFRcS34HwOSjZNEXu3FwHhrFomtRSLpL4B3b+Eyf2MSL1Hty5Zw4KXsT5icR4p3g
LYrNv7aJf5b6UP4hx5+XQ70U8i+I3rzXCGbOSt2UiVMat1mMVBFU+ujxwr/pu/3/M03xYcAehF36
KHQh+9QXHRhgBPPG/c30OS0H5CIi7tLb5XBmUf7/dEgU6Q8p5soHSGsCyhgk8Ld7SQNLTLewRKnf
P8lZ0Kh6Mja4c2B1gw7ofKSyxPeAWXLLPilvgM6SIpAMT9UEjroJinIlSgO2XMVSTsEtl4ebJs8J
G9EZnsHhfRM5v4W6rL2XioSySq4raKa83Ee7+v47igE+JTvhLmK5dDgq8fn+wjV5/pwHqUDQzqwH
BjmLWNRITg58pyz0jwONAYI5M2+1tcaMyNLk1bxbXq5vbqYmsaU6i41addufS0cLx/k4+TT26Es8
y0ugtRXpd2p81IdM7rF7g84fGzCCNp8XvcVRV8FhcMDuZkbzR8smvf0ZnPRjhYbWJIMmzfPB2rMr
81Y8Lh0kB4yCVw1MhwFoi+lHROhcNzNJYsPJayv9ZUWi7Pni08PDfixh0c03OivOVORVQHHI+nao
mOqG8itHw5ldSALpYslRxuF22QBVDZDj9nIXH7UrxySY5eer/no2kln2+O53txS58augZY5gJY/b
24zbRK9D1+MO4Lq+1kxjAWUMTusQJCJNd0zfpBn5cSyAFGmc6vbEXM1TaUBhECxebjqjgMAZzKsE
AFPJmb7hWf7bzQyNiZt95Nrl+gQ6qU406hsSb53TILvanwzVKOD1b2B8G6Wj3EYvBEysXFjGQ+vd
FcfscVMk2U0SRLyVJM46ma7sn4uOrtODDwZH9PjRuh3a7r0ooxucvFHycCXcQE4TKEtdn2scOUs3
JhtpL4WKFmEauvMGwOShm/6PeLKcXMrqAU+/TnpyrA853cXKlOigr6rGTHPzqzrss4WExX3rsGgW
qrvQ9aARuZDVWBt8PkrPUEcyx6unfKYqGv2irOgJ5QuWPq1Qx215uLBBCI+A3M3NZO7oE5iCAkSw
/sktc8jqiGvBH8JD8jkmEsnilD6cLPOOIF5ppDGTzmKaX/udz+4L1GygXA4HWMT8BvzUpYJ1FTza
Sk0ANcHrX0Gh3+Mt85gz25OBDwTYvvgGvsr8EW0apKZ/idXtxgzz9IOwvhyyp0U6lljd5MoMtFjg
NK4Iz53f6cEE47cQGFZCAdBNdwcToHR4mgVURzmomqy1m/ZXwa6DDn1v9tvVqAJrva1GA51PrhgI
3VgnwYBZlalzGoS9CdqwijGLSvqQkoOXlk5iB8x3SM5wPyvRF9e+/YdFSoV0RTUqGKuMvtJjdqa4
hMtBGKAmS4MlU78Y0vZ5AJWtkZhEoqQWnhl2t20HcOE07ZaazfYquNOiW/7SoAdj1sr7su30ZjHv
JYdPAkq904Rbk/F4Vkmpu0Sz8JG9bx1j2GXgAKdlbDgPLL8wigk8ipo5lf4vKjHhEeH9vykbCPsR
3GdykFNISk+2mb39v940lF4XyS3ApnpJxwhrDUVqf8A+Fhyp8SsDSN0w+3nrH0ig0jMt7q9I2NBA
g1D4V0XXEFO/uhUcIXF0eZhZy5r+DQtfeGcysQ3dw2QJMwFLBfXtle7fHXUEqi+5EP7azJAqwpdv
QOQm+s09oLvxlw+ADArqT+/mOkdVe5DnhiE+SVLmIwOpU9Jl8ghIUp0FKRvVgSaZ1UmgUxXJcZgv
Hjh2VII6ShDbkAe4raA9+fXp9EybEpTS+jdUEUqoAq/6cSCKpvnCquam54pGxopJUVJENWEYORjP
4qdWg59vOOnEPLF55Rcr1kpbMUEZ/aHljOt8YGh2nmR2ccnwr6xwB1TSsA0BaOSzmPuQuJ2qrcK4
Bij8X3sJSWceq41Xa6OpJANUfHi/R8BFxZcAtmYFo6DoaIAUKZDfkRQU5HbkT1M+OGThcLChVVAo
cqjBGC6u2IdqLtSZWRkK2y3XMGvD8e0wZPP3l8KWM1EaAlrpRakEdsFWHtLNSf8eDLgTV95uskhk
ZzYYsedp8YMBPKdH7hpy631y/AUwfCHw2H+LNYSAsztm/bSbFouTr1m5osFbb7xaUunQuSyZFRsp
zuuJfLK4r65Fm7HWX9SuLq98UZtW1kI6SONkTaOk6kKm3ouvj8OpBe/Igo6YM2ghWKP8n7bnqu3t
U87msUgh5Wyim1R9HbicW6v+0GHtPG/VYwwwhFFJC9qelfbwM3SClEdKN0E71xNSIZY8QySbu33q
HYZ9iS4W0nDmstCyDUBsIV12Iba2K3EXom3YNgdgo9ziS+wZULb1WczL4uoZW0MzDfbCFL0aHmSE
plTPAK76tJjFycTXMpGitEVSuAEjxCeNZyv46Uk1NBt0O5iyiQKyydC5ktgVj5/4AjfUWfXaIDaw
Fk/4p1Ot6hwh5MlEnG3DiP5Zzk6Twc1e830GptETARyjo/VEy8fm4ed5/LrshaHHHufs+8E2Fuj7
KjDhW+bKdQ2XgzuJHrqM7rnm2gWbbShGsa+6u2UYBm0x+OwKXQ+0/OMWg5Pqf2WRUEKPYWuOBYfT
iMzxZHvW/61/XHjmYz6bhfQUbn1Gb/mE71IhFRtAKTRwEukTZTK74yagYj6WXJGr/wu1x43KUWZ+
CXyJA9bKGarp/PgGsYyUEPNDznrC8XmsV3BVC0POpZkKgxPBvixwmkHcTmfthRI2IrByqe3GRq7m
LiXC4GXARiqbt1Y+VadCk+FGyz4q97tjae1ffPdL1S3lT0uFfkp61AWeMkLPRe07Ho9kYozjwg/a
jf8NZYmPYoAbOVpBLxDTX3K6OtJ6f6R816xbV7IfP12K5kpjqcwpGg17NTJ3dpEX6QtQIRlM2fv3
q7DniEZ6pTHVtRx9CwZuw/izcDOUtAkAy5eCQklQDaaOzzduq9Vg5RCFSJ+Oyk5dALRkfI3V5CDL
tCs6Q3X8ifNwlDPYkgrPZ9k6cIh0wlt2S15jShD6C1HngK+kgwXn9KfJoQxgPE9lsUzTNUdf/DAf
sSpF9gt7e2TiydFLgCiiUnbKwUCuNXV8Ah4zVrzWFBnNw6KwlvOwUXu9fNbXIN/Z6oiBPpaCcmAr
fAoC3Qz6y5ajGTSGMZdZr1FWeqhkdCLRuMfBMeDROQ24rv2PwPN0fXufzP/qdJUWmSriVgMNMfgb
5f0MyxeAP2NosnndwMpmCs3tiEcKeIdENSn02LkXZjp02w7LrAOOas3XnH/KyQQgC9/jWVxU7gTj
OOqRwIdMLY4qIyEngettPzzGiSOFmNznSWyE5LV9f33+JjPDSFxqSBDvl2lCMt2PHG/LaG+5NPSz
b02SZ1GrrkeQ8HA+gYi9uQsYRICj+4g1Dv1eB+dATsb+ohyKDh8EaDNN8aDUAhPgZX13mZF1ShWw
eyChau2YysqjlddnKKu2VaUjzieEtpXfHQiA0tNEpsajMDZaFAWWhz+DhOIYItN7HrBAByRDjbb0
GWj39dYUEy8Fz7mXNclWcvzTDUgj9rD6VQxLIh2Md55sKQrdVlU//EK3yi0YUwm6Q2kbFD+cWlhQ
YNHdVRUPAoWPKyWuAV1tsunmth0ECeYcdqcKXDeWgltHlViXMdRSlfRvPrafCPxcC/JRduwWRqnW
y8Rltzk6CaPbtg+ILA6/8xdaNlI9/TlG7nUtg7mftKkAGJb3ytthFxFhZRxAHemJLjLVNg1PvE8k
l6a8mY6C4CGnt2v+g2ZUsLQUygxjyiyiGIEzT7WGdMRlur/53Fim8r2MN4mGI6NVXMQaHa/EuXyR
LOO3rK1pmd+jHHcR1afDp66Q2bC+xYoU7GELOMtfICWP2vsIzdsBZ287c0F5UpnDKax6HKfo5TkQ
06vYMaRC6rXJ1gAQQMZdFyTOsHZZREtfFeHUWVlBTJ8chnZff1FbKp4AiObmiPbGNoH5BtLDNkol
8YEcmWnHV/0IMNz3Pslf+IvzF1AnK1HrVdZAzYrmE4MTh+NnQsRC7MaWFqrvYl2fsktHM6Fz3Hdw
+Y6CtLOLbHKX+5ZU4QBWFl3MRbk++CNueSJcidk75PE01dXKPU1R9uZw5+nWWqXLW9laRwBCqzGy
j/sY61z/O2rD5Z7IGQjQvtwDkxFTeIOl5h85E5Zo+J8NSIPtHns8ArwKxCgiEswJrc3TfEyXOFgM
iLjJN3rr5dzAksFySDMVUun976RvmxYeSrJ5ZuGQlFBXBYfUFUza3+eiU/Q6t7VuOnAbGn6w2sxw
ByfW/C+yspKig/nA6pUktBc52IeSAs5QtVzomBuLKMCAXAOIFqR696PFuAsWozK8IJ9iCj5E4DMA
+pDr1XYwy0eK1VfGWvpuIir9MR0zc8XfHt44h1vrLpTccm8eIxbx7X0NryueZpNmJTRhKjc7YwDn
te0+Cf5wTBqby4daPi3cv2pZx4XaPw1urrdYBYoq+1EXhps49vd+JmjOdKLkh2QwESBu3nDBMjqo
Faa1YK9STZL6YY65V5TlY5cexLD1FTPVpb0tOvRhsXIDJ10409Syo8EOcJBm3ZZWwwrB51Az6elw
twntS+Z1pdwI9QZ1mLiUq8u1moXuurcRD1laLf3jcwybnUsrHGKMQ5g5kvc/vXTkD7Q53WRxDtpm
lQ9CQQx5FmxDjUA3BxoEVEYzyQIaOTFdEoMpAGq5zqmG06r5K17ZaRYicvFKTxXrdKrfr1nS3SD2
28Q7O81m4deOT1uNe9K+uN7yKXWAXUrrCWrLAjytMEFF79mHm//L6BKew8hHdpbmGRHi5/908rTf
Fok3Wise75J44q9ksu+eniX8rYcABa1Bzue2uOjcvnsldyeN3eSTtthenlc2aAB+btARGznblM7Y
EikAO0VUgSqlihojHbSMOM1kjsZV1nfAizboBBvOO5iutDJZXpZYucJc8nfy5D3dk7LiQ2giACzB
tl5CJ+YtjNj9/0sF85Xi92855XUPa1O7B4bnYJ0lNXqQIcl4vt81WaVccpJnPYZmcXYkLFWAc9uT
RzMKqZoCRphtgQOLWXCJBDNdals1Hx3PysItY6BXDQ1h7GqgxhEfkjGPyCTIanUlFFs/W+8wVJ9W
/uNzhLkwIR3keLa4IOAjdMpi9Gihq3UT7Ulf+SdPBvr4NPByDgi66UC6PuYzlkUDqJN6I9JOYvrR
/tRIU4iHVX/6adorMJPwk87ir2LTXRMWAxwvLJ+bx4h7SyokEy3rfh7DMfu7iivPEenkD2i4yUMO
wP3Sr67IN5zfsZ3589ZXkfGn0+sY6/YxuUAPadxhTCeoQLoObzZfUyKK17SmhEFcb7QimBWvx6RO
snfL00NbVPdv//1QhKhU9pJECMj3r/XjCBhGN1HRAC8QVfuNlG1Kt+Pt7ufatSm/AH0ZD1zHVT/i
1seu+d43kZj+M9UR2p6fYEDOA5kAIqwwCBlSa8xLSCCvVwGSgt71Ujq6qM1N7PMO/Cx6XWYFAMgZ
ymCN0a0tjpSvGAXQ8XjbmTHC1ori1tIZBx/NJ0QWhH99NWDqo3wu51mLL42EIuwrLRUXCHZtgQOI
QbfHFWONApOG57GG1Qdl/u0t/CbInkK5mlCNTOJZA0K5b45v2eF6imLvmi7H4fM3pEY6kfU31JaK
10/pSTiqhmACUPWFsuTqqy6DJSGqXU+D9Dq1wNfP24g665f2kV7vBALUAyQ3Mb4DFHf+nnZPg/vW
h2tzUrIa97Y6bCfVxADZqsOzA/jK7GszjIR9xrBP4qCJBbE2pptXHKi+gSTd246cE8ONOc76fbC2
MGdvNbBd+72SUHrn8/OR0co4xAIFD0kwsrhTMPf/6EJT01EsqJvpwyzypD7LihoXXr/vaIYyo8BZ
zIxJ2qjz/Gdwoh0OKxSQKTXBsrrDD9DpOeWzQGdCrxAbT0r9U5zjmWiLyN80w6ux9JjTLMYPp4t0
OrQz4dpSeHzRJhTb8mSAyTeOSCRPNYaKI8ftjOxHX50i9AnPJ92H7DKD41rgkI41pIyqyCJAqeed
Nbf6liFp1Zgs46AfuJN1lQdWQOkVT979RV8INEF5pxWkWOVRF+2pXook90rRYkSwnYBBiAxluOJE
Ke2I23YfkuxpyJADJ7SYYJGCZ4shzoiIeNY5ezI9gBSHLK43O1jJ2Cq9iCvgUy5CAJ5qQ6/5Lrvo
x8N0XSviiw5jQ0Ez/CQQLvRtkSKoyPbzeGiuWP0u/tdCuFhHvqmYiVqvyfI9HFYUnrnZHKeV9awx
OoIpXOIkQVZL5tQ3mBB5qzWzQh7gE3XpVRNNB6wsf7oNJX3JeaY84Kd1dcT/9B8CoUV0AVKAdBWx
pqv12c2CmJnRiCObL0RKRHg+0E6ILreSSBfE6KzXwvFEWg5CzyDa+iAUDjfeaKEsd2LSlewkOqnT
0PNR/t3hhDV2FdTj22cw47N+Fu1MLiMop0EftyL8IbpCB6Vrw0l2vmjZ+S6nwSfI11lU7rskJ4x0
XO82qen/9Af/pjP3UjxJEKKNwB00T/NLv3UX4M7e6GyVD/b4MFOCyhTrUauq2JTjMQEYUX1+zZQ2
sffzQrx10JOBd4BsbZ6LxtEdKTye3IUpyZatBcrLhJsOCp32QYJWkADTYUrdENwPFRG+5dtSWxgC
pxuWlIarbIcsYah91VfFDEuAwZVTFroBAGD6ZYKZgxVbQRWU7pl3tuK3xzX4uJHRR8YD6w3sagHs
cWoto0J/CtgkZa3Tce+5ATRKg2Ylwjh4wQ2rusFCHdw59fivTNovwicEyCWeVI97t+dYtJzO27PR
UbZwqY6Mz1CwjM49X3Dn+f0fGeR4DVYxDYui3+TOJcJWrmlc+sQ67dnMhb483//MUj3zotvSssjH
fDynSzEfDtkBon437Rd7Qq/MXUGjmyyt0tyilTytGna6SCiAF748QpE+LWUBE8Oq10CLj0wqfA1+
ADWBqsXEboOgnKydwRQZ4YXGvQBQzSS3CvnuIj2fvfOsm0GhnG1Z//MlxkTU/IVGl6ijdH48fVH8
5HeXvTKvYK2tJXdsffZnaQIeV2eSyWQ9h01h22RMqiT6VletZIiHc/E7YJwHyeCVT4LHvqY1106y
H7TAfUU6EEHQTG5p+92eskIhIMpPmr3hzOrm2XiwDp5c8qK1CoEw/Kqd7BqsHezUr67OE9ZJ/Tio
d8bDUwrgKCDzaKrpg/6Nq0c/E0p7+q0z1FbQzDjaEr6hZCbA/B18V8R/5gY8Te0zjEMbI416nt7p
dK5zHuSMb4NeePNmhMWpgH9nUsPfz6Mof4oOHiJBzufonqp+bqUOdRPrCrSTbr3Jvja/LCDD86vL
2qZw0hgAIqS0nzhNoNCNuEYlXTYmRoZq5JKvP6dqoQVV+ntIrfgG2C7t1RIdWyLfTJDX07VH7yG0
XRFSMWNf/zHmozecwl7DBghEW4YMEGQMcnVbEjHrWI1dK0vAwzDeMb6GB0qbP54hbzQ7byHSb9NA
JiGAWZ6HUPpM4Fx89eLeVrCvvSEUHtXjWzOyLNW8q0Lv3VDhfVArT3qhsmk7e6SXUP9Zw/qpjBGf
ty4e36No70yM7zPAMYkDgnGyksQ47CrcrexG6WYnLQgdIMPx+SnX4Fnuhjx3m9hxg7SsWpJVk0Gn
WvJQU9lWjSuhvxsQNzVKoBjNnRHMkL/QmAyWAJdWq1Hncmnvxy0D1m1vdoENZnrYfg6X7kfGTvpG
tw8+dsjR5prazb7cGXETHWVaAgopZXCHvSkj2eiNS+bhDBR88xOZCeZKMnJAvj59+GLHBUAmwiGj
GRI1MMhxKyoMwwDNADFNiXSkqTIzk63QkIQN6nrUBLfZMlqOTShb0G9BopY7/ymQmv4/uKl3AuJg
g/cTFb6sokcLXpgR7VWeJQvH7aeZ6Z7gaD4yrr3HB+xrW7SMQs+ljd4ulWd1650odB8Pe+hnX5Gf
R1yOlDJ8H+1DV+LaeK/9bpCQjrIb21tb9UMoeplW5xuS2lB58NBbJnzRMGZ0WRPk6fxUvbBxNpjs
BvMgcv+srRuSvSH9t+HMbn72QZ5SxVlG5XG6Z7XPKNg0k0lMHogI8TBqnRucCzfk/pgXQAtn1DQI
L7ZQwSdXzaMxfTjviq4eFcwzkaJXpZHTnTlfVSWcJuyLSiWTNfqvYvlRCg4MvReYCAr1sUuT6LTi
ShRu5/PO6+UtnbkrWN+RdkJobNc8o1TRMMZku6B7I9PypsiKxRwj+0B2/HnV+wILh/meW957wVU3
Tl445kaHnFyqPvXLQesv306BCeIokomF2ci1mHP0flZuDBISE0jARfBI9XP8zNOItT6VBwOcafyl
hg0xhqTW2h3cvSdMQrWJvkK2IEoTeLv3KehI3OOn79sfMsbf2LSzIBIcThMicNWMHupadaADG5eL
TcaMwJnGoYTh3PPOn/WOB5U0OgYzQe1BYlcCCe9nEPfk90uWhIvoDlvL76DitOxtaRK48ko8TmLy
WldnwzL9e83jNwLnNYnJzdXf22h3nOuGbTr4O8rF+0Q4M4bb7yfHT0Ok/ov2YrNzmT9Q1lanbRVv
k7/2e2sTUGSzUrTj/z0kkQMvunRJ9ovFnxibQ4cBa6t9fRLXsP8PW7MyR1g/laWeZOqhqW129Lic
o+DirFC29x1KvStpre7EDdhhPkTjn/e4FJvnOUzxRw0PqoaGcVaVTSptLfRgAOvRRGllH90Mr2Ab
IieIqZYLzHQQNzhp98CGr7bCekfxp4KtU6JU54sWKkeFqg64WXYE3dXggEqJ+33CReILzHDdj2CA
3exXo1xRQexSCq8vfZfOIXXgTJb/iA5vG1bdy7k2tClUdVopGEbw3gV9p871BgH8zVZZp5lDElTK
J9euJDlnzpoMUl2WSIzD3lbRdX54UQ0nEem26IgbxGtiUkE0/VxB0PXDAtIMr1R1mo7vQ5iicqui
9VhsEcjzqQHluN4TIAD+4XU0NTFjBqi9AFRe2yf+Dv4Mt5q+tcv7hQv6peLtk0A0+OZo1jWFI8MG
a7Vh38bRGotPzc4sy/jsoUiMOOyZUjpgx2QE+JcMcjaQf01uEr6db1r/jITQjk9uIn2NOMOG0F8z
Yl2jEua5RJtL1j7J0wTO+WNt4CKex0YmduYnmx/vHQK3llDAwy9oGZ8rq94xzCh91/biXqrekAnm
yGMWssMqcBz2OMaKqPTSVHBPqxVc5mxsnJfM0fJkQwBea8ichmb96LQUPHLPzQmYvmPpM0VirMQX
sMHOSPcCK0KV/8by/rdy/wWuHJK4OKTe25JuXGFpa8d1CcXGN8bjXxHnX49aIelnIjhutiN+iiHh
vLsB5FvfFldGpXeIXWpWqYbod+jbILGVHSc/5NKaLRkTqkiGgbWf/KGJbFgKbf10lS9VEzTkt/Xv
88b2pdOybLlKwgTEPVhousU6wovDR92BRC8Dn0c7DhxcFgMzSlPjGzmOu/GqL2H/ETyJoFy6LdQ6
n/44lYFhstvIMScJsCL1142dC2AbfGjpi9oI0lEfADZmjxqSa3l9ofPnwxAqgKvIULkFI4nGR2Ld
fnqZEqVeva7WrRMWWMcw4s3n375f50nKWfPJP7N7zXpCni8/NrFPKzVRiI1RyV1uys6JXCMD9ZCT
msWKavn3Wpj5PMil8fqgM5xEIddUerzw1S/WvY8J2FwculAGFtbtlfunfLH9jROd/LVi3i6+vwuG
sDw/J/4hMAQANBcCjf0cJNc2q1vI28QGYcNMFi3AvMhZ4N12IbrmKVXcHgyXVVYohqNiHcCMvgby
4tgSf8ZhrUqMzPzxLQbmmoXcecxToWPv+qUPZlHKpWbbdzKNYmZEr18UhIfIvAt9z8tTi52x5p7u
DC94jiRrJQlpyCxPzgws8rO+pYE+ADS4RvNgqf7Rv3fJhn9lmXqMCS/9sGFmCAvWrnZmKhhCdna1
yILa8i5EgzAMrsCSJD2LQ/L/+8xdvb8T2im/oTErCEfvBylXc+u6ggfCYVyMbkbfyMk8+BZTag48
tNOHKpVbXucdLQqF55FvV55MXouC/kP6ECSfmxdSPTmEg376HzHjW7FQvvU5inF3caqPYBaEYfZu
BkXpgOcs/FM/6174HUAk0klvwdGgQtG8HtJSWyoSjbRnnRlw5mCSdc9ZVItGce+QaPeeVsx6Uvmv
YxD3QFCKvQKh6Na25P0uD5usNBn9X2RuKiInLTykJwR6xkvdD5ezuTAOsYikE4PVzORnLKgnI3PQ
8e98ar/ZOnODhl9M2NJKiSzHuX5RyHY7sQ1z/osIFfab/HI3Lt1uaOovCNov/issE4Ey4DL0J4WM
YF3Fksx2UZ/M45UPV0QhFN1LTfJ27/8Nl079d/vxbUFsY0rdlfrpmiLjIHV39kgngp1yCNVP2iM9
PsvEhWD5cjLyaPVAGg7T5cHl5zzFq/Z5uVKbPfaF1VZusMLo1ToWfzSdfA8+kZxjieLMhaqAeXBd
KlHbtj9VqO3RkgYXCk5CK1o8BKh68tiInjb1JZLV7dcnBf9mP84ZKTLUIYrwCQQ/H9mPfOMdcwAw
DLQ1DKoupmW5g8rzNBMpx2N5NDXBDBUPIndLZnxWtTfUpuGnKLPn5NmxZR1kHnDWHSYef4jX5oJj
bYksTVblPS3CHJ5q8Rz5St2JybFusgx4Qizdi8w01Lu8x/BZwURcmTI93NHY7/GoplmPJ9sR5T85
QQ2YddB2EKT9Do6vbnmCeiK/Uv/EsfQr8YqGis8wnWhW5YVGs6n2O5IypkNENjUV+vyOZZQmaK60
2Tj55pXvjqzKyXEASOtkJMSREf4QG9B1OrHkA3RgK0J4h7JcA3syl/6MoUEeYZML5lph8mAwqiUr
o7AlQFWkbKgIY2DZwZjAL7XvjRloFsgaC02R8+qhVD6fpD/YjEhMEHT5GXtky2ctsYfNVgQ0ozXN
R5JArIsy2XiVpY5RWQINIsrjKwQnapj6QpFCP3uiuZ4H6+r9oT8FsusTixkm7aB4jlfmm6tq+U9f
7naJ0zHKRHEOKcwnH8BGuSw2H5KzdHnsCFdnmz50JkARdeOC8LjcVn2F3emd8W4fj2TGwTwACoZY
geFJw02H1VBBZXXfyxkvK3nZtjSGh97ATDUn7lY/WqX9Q0wL6BksIRHNUA4wSlWd4+UKLvJkRa3C
oiFXWydeh+S8Vpd81WGF54Jt3BGRWE4GMZpONkCwt/l0A/VthpQ7BtOWpvuWmJdfpLpB3wnsdXGu
mL46yIyiG6wFY6CwPM+JrqtaLNpuqcdk71RagzmLLe8EsgDJY2QZIEgFDcF4eQLINyRlxK/aOOQd
wZlTe3U5UO21MY8P0rLH7V3nyQD6ivvMAnOxovCniQXwe1yUFir1wlZYpUj7/A6zIt4fgEPDwGpn
OKflhM7drwXzRQKJ2wtGqPDFj84KRPNie3hKzABJXMdb7D51ZuLKmuaCmvE3hoat/C25MI5dep96
uT+SFzXesQ85jkksJJd++z/GQD2fmdJ3StIRLSw6kAbB182lMg3cUPj7NG+Jt+8XzM9PxpRd1f8V
RscIwNfoWqxbfVy3xhEMHNVh8Kg82OT448+bNkLyxZhQmBi9kI3IojCB9KmBveyEwsXknuZKbzxE
X0JE4jHj9vQ2VAcyyZjuU1WumOudwuNZd+s1VUtiw8oDicGaNzJeOMkaYoChjGGDCVuUg11cblVz
qlOU9ZD5sqF5y6lrAjkXx/0uaW67xYa6Ri8GlB4JuIaaSjVbYvfJy2PBNhJQ3VeGtal7IbXhhCgQ
Gx/WaeC257Dvsizrvp4Ca7BDeoIt4ptsA8HKIFIN6gatpQNhPtXzwUHdTirbp3/FNFQhSvxJGlq0
RI4zCCZOnBsaY6qX26rqPy4UqtSsHMTk62in7mO1KLyb1UeLmcqVH1I56Z+86J6r020IwXfSBCfu
YFZ2xQLjTijvaY9vqpbr+gMbbOmY4YtALpvxxQKmfCT2KYCNttGXFMYcB5bbLCyU0rVkOmLqiviF
qnABN/18qGuFjewkU79JVnvLJN2hiEdOxxUJzAZ0xoOXIWa0OqON5i0pmc8VstSIIFX/gwrxupKa
37O0C1GQxFnoTMSzh4Eun3kD+XlAVhuiJNNbXAu8/kz3NLD68r1le3AtpoJSxWdZJA20WWVzvUKW
AmuJoconB2rjE8rzIyGvi2WYeKksH3PRbm/Cp7PcH95xgqZcH7r5+W8kjxRzIhHhJxgJN24PUdEp
bTHpA8J0HOsWHMElUs/UiYr1nJ5BnJxn36RWWdjdoz1dBZdpepdGSJRhi/8+sHcY66l+W3KyU74H
l8KwqB8rQztFtkktTTgDsThdeXZYjIKG8m7ivyKixsUMw9Lmfy2TgZHRpp1Nsnq9+45gZCAwNjDM
fKvXL8/Oxg4tLyLN4f0ts4MZS4+0KjaMBLWNpsabGVQM/MTXQHQ3iNPipanwo4LgD02FwCesBPmq
tbrCwsGwBk5U0MzkioP0BUL9y6FgaTZxRMFW2luDQh01TMnQHD6QJR/6OvkDNJIvYOTPqXax9G8O
QQyMemPxHKEg8+X4BvwxalDcY0pHR5aBzk9tm5J29f2IY6V3r9B/K4ee9KDW5ksEGTqGK66fJURg
ez9W47TlCjZVIB+gtMHAxlkWKu3zUuqnRe49YNrXX4HtRzi6tZFEm0mv433W/CmZh6REnRrR51Ma
PkQasOlAbsvk5TYlOr40PBUkPUGlwjsD5MV+wDdbgthGXSIZZ8tIsXLPNthoQCnO4vCr1ddIyhES
JQcc//AWStpHDpuapu8Tsu2RyLPP7uZ+WUzbd3XpTWdnSTfrK0JvVdtvRBD2mrYchrz+dkDhL7Qo
thJnZIUAf+whmph4tVQmVug2to6oyVpFcIy5ESvdXLFMWk7vckutwxjo2a89Vj4eUIsHn9ZqLMCg
8GXkWYv7INQNLHgtrsV95buAcR1/rQtqmJMPLXHTFkosCKNZ1b+ZhpHymrNikIrcDuKKOT8RzUno
YSmL1mh4qS5gKt9EO3v5V0XrF8o9iLoTA5a0t1Xc5igI8JRdxAFApK40qCh4A0jFdWlwOHOT4tef
5isaintVnFnC6/CUGHRwEDg9vJRvjIzBailnqTWVFdbP6q5kBnucqJpF9NnPbwyq/seADCgximSL
DSzOSrhQMBPp7pklkOoJKibKJsQ1bYTGhnrYxPx2YsUKfP1DvUp6tsIalupEXhUZrpfxYKgeQnUz
Ai13qiguQkX0BdTPhTCbw601CLtpiQ7xz+XWIE6zGMwAy7dmEir+pdfnzyyUDs4rTWcJpUjYvasp
c7HiSPaeP84b9+reZKFLwPfZ7gN5YBK8BXYJgVTFwP5l8l5gxtVYPoL8ZsCm5xx+Q5egZykpDVe6
EKZHZDQ8fJRLv3ekdJiisyX6sc4VqRa7TysGW0azzrHVT+WoGa7xj6CKW1Hs2Ifpg247jL5DPssz
fIDUrkBV2vuuB5doV3sIVKZ3JIyfWrLmAlCToFfkGOJ/y9kRMZ7U62hqAZboEsvtiXZgAavp2Tjg
c1D6T6SefNa2gXKeAqprJX43z2Zgct39OU1aQzz2b/Pnkg3Jz1zSiNBhCGhANBoEQaEbedsrQVRd
3J6t9M3JwIp78I/64eXth79O2ZMwH1peUC4eJ47IJ9EIILFo3kiiFGV3eU7j+RZXJ9J++ZA+wvdx
ze6zBpvaoznHYPmqpNS1LbZMd6bfxEywF8l3WS/y2kh2vzr0qQfr+0XVj2IGfcglrMVjgL3EwxpM
2WZsfvo69rb/FWGOnevqLXf2DMp8b4J2qAbHyKNbFrh4gfEjbW+jCH65Wh8TvYbFbuYG+44Ms/OI
/UGC4H4PW5fb89dIQnOSJcVgnt+i8paeHWRXj1YL6K8Fai2jco5F16HifY9i6Q+9w9qx2obYmbaO
2SIXKP/GxygKq8lD+wq1FvjstpBu32xKSvlBDZHIOh208rG0Nq4eiHWmUfAKN6hHh/DtpQfWnOT5
4tPWPIAkbFInXZGK4FSHaHapPpA51HMLxEHa4IRmTYWAdLkgLAU0KUcNDkPm+QfVwIMuKGGv7guX
vM3al/EQubVKqngeNRe8JzwtKINZs2JOLLEjVGj9sh9M3IV2qQptfmLP4ScAMCA89N+l/HEWAetz
9/lSElisYCGjBylP8ehf1RBG3MPsfs1DngvDjuNqnr08VXdYjOmJDeu/Ei/bawlEGBkaLAVhHLTD
r171UBnddgPF5MeZd5vB/L0tE43hrm+tUCUdt0Qs6rfwPeCm+l6Y92k1Ox3aDQhr4mhssD6i+5aJ
6l5OSHTm2bt9aIl6swaBOcKU2VzGPJTcQdKIEdKEbrfQlpn7IxI/UVGoD/occFSF3kE/SUBKvdsZ
l/KeAIkJstMEz/RCezp0D2SAZwQ1AXdDo5vc/D/PwCpmH2RALNyA0YOgsJCBhK1/ABX/8NTSXhgy
5YWIJ3Yqd7orkJkb3jboC1XRGRm70nM35bI2QKSw20/Tf6FpmH5itUefsAUAaMvfREg78Tq77TmS
Td/Xf1TXlevkL/pe6KxFlF5PMXcidEyXG28nBOBuRW4rfIeq+CZEtLtRQZo76L1FMONT3SUFrJR0
uuS1BVX8oEmCbSi0XBTPQbs48slLQraBTen4atPGo9V1bau6vOvpdefM1+4GHwj773Ef972Iaykr
yrWLOZ+cBsl9i4EYoUoEkVhbkUDl8mSE4/3r3D1mhct7xcoY8u9XSClV6T2fLlyrcRcewuZejXAy
ivu3H0IXPxqSofEfpZdpQWnQIyA2nxSTZIj6uua/qjUVclGNZvhkXsnvn4lAYqFHjmkQUu6U1kny
ZuFC5JVAXcJdKDhCkWHzQMAGT8JOOYo5WHQitR0dotToIOoYx5ayNx9KAb8vEKNR4wbpJk1UbLyF
KQugrqmfm2+ynBX+FzpMrBn8rUs+7B3ZlH+kJc5fh9I0rbQ7Xq+xB9D9GkGQU82g4cFItemo8qxq
1Owkqq1f632kcrJM46SE1qVY8PD4BaTXk+MxTpwaZJ+ojFR/LhXy//nb661F/e3YGmolNwHKWAzH
zr+3rRU7eiBl4wav5Yiy/vZ690cD8RsDA6cjsOLNmicduBbmf8y4CCvumPYIbLxe/bY25S1jQXbv
7nQ+ywgA65vmy9XSKUUTAefWQaemobyRlEl++ByLs/GILzdnTHioymk+I5V00fZE1GQTNI+2/McG
Tl2OJdXuN4aOcGfZyY8VhSbT8sDI2ZxL5kKyThA2p6Cx0dS9qzGJDWtVA+2qgMe9cnFlbJ+H83dz
yPFzFEsvg/VV1WplYnCybUoqX95QkQYj5jJJZ0SZdZdxmDyK2Jlc80D42N9g4x9l3xJfL8BHe671
vvLryNF6j9rKWz+gcMogP5SbUF3JSEW68yo8amSs5kIyxbwHU3wmPFo/ZpXkCLwGusJRpYFsZcxB
FW8BxeJwvYJl+vPwIiaMbixPwJe7YGmmR2fzm0fxeKXFjO9DKVUo0q5HeaveiX1MjGPciagg7Bxl
KTAePoUXJbxPQVaQmyHn6CN8JDWK3Adt43AkX53+g4NoOn2x/0ec3YKMwqvqWMU2RRpbw8a77erA
wMHrAZy83yjPM0qP2+OEWDzev8EM2Vwn6/cerRHUJKufgO9/ldzgSc3fkH65w9ZtFaktCNdpmaNK
kDr24PLMPZoW+bcHJEoFQBWqQpgjY8rio1z22V3yqS1L3cXS7/J2zynpg7dkTGHzevhzUIZDFe/F
lMM4kaS8iHjGzcQt7pkvPugdJ9GKd8mCpUWPhoi5mEfZaRuedj61TIBG3GeRL3A9ROt7QRCNQpy0
ug6K3JsxtnyUNYxwLJTOXQ4v4hc+mJF7J4ZtYs/bFMfcMieU9GZ9vL//Fc+EUnXSEfwRSz7vQUOb
aPwC9It8hDsVPnE/fbSzK9zk
`pragma protect end_protected

