`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
1+GJcjqb2xNweLV8yg5GWXgj8dCDk+t9Qxs5RYzJy51YunIs9xR9knZjn/Rx5sfQYK2Xnl3kha3I
bRIzpP7QdEp1WbbhMxhm789Uy1b/b9RNRkQVetgGtru7rPDKYrulZpNdWBYkdLhrM24P2Q5rA09r
UZGgi8S3Et43S+TAMtoPxcxDZt/4jPv5A4zyIqRnlSZZrvXnMFZ7yTRh60rvjwt17RC1hFUZ1n/c
LSZmWCReJJhzshMlE1z4OYt291z4vuaNKYyMNm1Wl8EO+SsB5xPb6OmKnmB+d3AMMacXeoKjv2sz
F0yJ8geERx2bcJCGPhDlEAJgsTvO2eL8XRqiHA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
ue+5QtFmV/7HCM0xNCsVG7tBsMeDgeDGY5WcgOW0ZKnVAgDmykg7o0YYsCtiV2UVz0txCiRcz/BV
heaKI6ZnG4CIoWQab2MZxAI0vjOvt+z6TpYSklwLqMf0V877PmxpyHzIBCGqy3sxONuOFBXGQoAY
zo2C+w/S4iBgWh56NtJj6vzICkhjwoxsoNEwMZoSeOochpP5pcu3XeV5caGsbrn5dbvWsbYF41v0
5/nvJqMT5S6jaROMe5xBrN3fAfvUxq3MupKTQMKW186o8bZgQBe1bIj6z5JCsNzhvbfpToPI+HvQ
5cWkw3AVd2yEDaZBGetq9vAXukXvYCBCV/XtqwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
DK20HCzOQTlN+05tKCWSBvRqcM2QDVNRLNLiIWW0m9x5EJb4DbSqLw5AoeqUWQvbakC6IKy7YaKh
4MBzSH5+GQ==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NVNw4igxMe9g0oqqcYK0tQXu93OvDI0uYulSfEfkgNL7Y3IZKoG3U08cbPJZ08+LQZYW2OnZnAPj
C8BGEOey8cUhznw/EdmN9coEqkw5PAt6d5oTpo8q+ydzuN1WU9Z6t/d4k/SecsDXcx9QIYdmlDVO
/porfO0TibY7JVigsIJI+FqjswbZ/cbnexA8lRGxeGCTGfhtQayC25/GPcnUKvgoJgPdTg1KUEag
PRw8doFCOOdUgi1z5FIbcUEX8GqyzC9Je8rDfSQ3jRYRh+eFgvVfoJjZveqGvp9wJ9DIAigzqTwq
2he72MW3KK/BDZA2vp6wMXEAyX7Kd7xqTY1F9g==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
pVQxd6m7DOmqSkkiZ0vpEVfSHnAifK+YzE2+wynBh3WuajmLioPnJ/UcuTzlQAJACvOrxntIdZgX
f8ZosbZ+487aFa+5cKLYiPSqpVK6mzU3ZgjP9Qe+nB9P0zuKitDx7BdCYViPxCp5Yuy+3kL2s25w
zaWPieOY+1UyvW03C1KozJJXtMmV1+amVjA8KG0Z3/Ot4bm92ScFF0savWKVBaq/SsklNbbDMaH4
KgsjQqwvMLSvsKQafiOnSQjFhd/1C94vlBkKtsjjem5BY4P3rEpXGbFbjLUhw0PVZX8Dctf8xYKZ
xCagGH80RCan88ZutTu2ltUou3r/35VXshPtaQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ICkd/mEcZbG/At+2ZoYnU7qwtdSzyLvCWxJnemhqGGwKARbIAHgNd/FFwEpGlCU6BSth8MMJ2+pn
1P3piOBqaeHsrNgw4dJBGqaxJrxVX9K3LoOZo4v9sRS7QEtXySers2qZXzCsdDsdRPNPsF579ODi
Q75tLU7fO3LTwuMA0Ao=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Io4j09GZku7TvxyibhDSWm884OfKcrk2NGSr2KM+GeH3fZVvSOiPvHSdP9pFALpZ74Gl24/PB2/f
MMcmwhuFANx7PbFPuO0jigoAFHAsDPR0cD4d/yHwTslWQ3aHSdWbxFMgJT7A0NQs/9cNXs3OdWI+
Bx51932SgduVO9EqPpTJ2cf80DFdFIXJNYdJZtxpWW7uz71swlxI31C8KzafeD5qS6vlo9hwmd1s
EErEbX5Dukg1WC913kRbEnm+bBUmsTYQtCGLHq0nGFG8eyVw/ROoAT7xg/9mh9DXy88/eY/CwAX7
KoWtJbFrFFoETg3Cnrfl4oPCrEK02XAjiyU0gw==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
GoOkFPIU8v/xSW79tGQrqczaUSFW3//Qi+D0m/SKGl7tmX7V/QfyNVa/dDZulSNnZreOnZVulIDR
sf+qHMtCyCeMtpNXMZ2v8FVk6obepqwrh6w94r4+10yKsy/7GSi9bSeXe/HfY45eBoOMCfu+ahaK
20MLZ0qMCoYHTbwlXMO5/hYiBmA7AImMVT3HwN8lD00/4XCcxemSNZWfGwihGtY7gTTee0ZQGR5N
Y0wxwykhmmIBIXit0ibA8SqwqWfr0rQEpE/Vj+ZHQAz4os1NhxtOmI1zHA4HisRUW5b4VkC4fmyi
cFgifdS4amZxi27p8LN0ygoSwVMl7NlVi6DrVw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nEAJZVr5NEWk/8uw/E5MHPdL4WN9Nqu3Qh46OWCx7ezkCRCBkKH+WHp8nJRwkd7vBOyGtcLKkKxz
zx/qTjzvjNg0OK8zJQlMAz+OivWID5IM+NQVgHag4XvkP9kOnkb58SyYwDmvFDGZ5WPoU2F+94li
UTHEBCbFX0093FLbL58=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KY2DjKqtQZqZgvL3k3cC4obeiEtjCwFLnNNI6QjUnPeA53aDq2UvfTcEj5CQrgF+yZMfHoQvQ+SK
3nt+MDgNc6kCav/7tW2yp9cCYUxkEVrYsemIGZkxFWqiMarbuf+6nalT+t2vrjnNgXZ+DXT8tSN8
Y/v4nkasYWatE3X9Iu+CCzSWzxQC+SpOZAPWPf0KwU5hgmvHPXDYP9e7Z87xT8DXUNw+rbE/5LSn
kpvOeAbv5/kNUNnRRQcooY1LOtn1XPj6TyRLgaJnSLqj7k+CDGYywwF3mcGtSu7AlwtTUDdwfUUB
abBQVOdjHJdGVDVdqa5BH7jq02uLaWiAwGJm0Q==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2784)
`pragma protect data_block
gl/PsdsUt+cjMOgz6HFkQJJFlOBmaFmzrBhKZQfXEM/UgoIumFwYgs/B0lhD3aV/JjZDnVv4Yz3i
XuvnOx8aP1NSU3/EWhs94eEl5ud5/P+9n2OUIZ0GJ1+xs674IaJ+Fok0kkTzvggiYXWskJmFdcDM
q2nF5B0J3TN8bfz2hx7jIO7ooQIuX2Nhl7Jqq0xHNbEix8eq+freDu7+rRHNFwHmr/0N901yMPql
Z/6OLJDEf6ozqSOudOZE4HnQWqUE9DQr65cAkokcjvGuzVhCUN+hGYVE3512WgMtTz1/bg+ozp9A
qNUs9N+yhQuLE4vtrQrar3vU2lsoZglANS2WaFm7oK5KBOitShWbi4AwPhPce3ZI8vS5nwfM1ydS
2XfVsR0TAIAkFpFqiwnDvJqekktuRY+ociDql4c5bGTXh3lRAXMf6Em/RwephTz/2E84Le7sWTSE
Zqo9JC8qOytDxm/UGeYNnRdiXJy5v/gvF6TKvf73BL+ubsDoBz6Pd/tTaarwvNBXS7ekbJWOO5T6
sSNR5OO6j1ubZrMVI51F4Gv9NxFUxJ2rKlmoI5jAx6oDATDFiUceRIplzcMuO0jVlfq1g9WVB4P8
Gx9krNAbJVA2BJ1jTQ1/Bk+Xm2I6BRvM0tNdZ/JiPZVBpxVftTM+gIQ99c/o2fmqvpJ23LCEltjF
gZyg0m0E6UBtsrvU9ua58JRI3jNmTUMYYXOFYYL+qMZo8mTCN/fJDye8B5o5NJ/3vEDOvWQeHb7s
lCidwqigCDB2O5vST6xwvGMAKVbRq+pw+uY/untf94pUrjSS0HN1b9Syv95Q6NOdun1dY7tEUJru
PzsGcQnLZJx4GHM3Kun9hdJc2zhLGpzYiowbrErbKxJ+ZltqFJ1S3MsH7eUJsZ+JoRA4MkWWEc5S
CE7W6A+0NRGpoXwx79GqEsrHk5a2KxlaOd/aFMmMHjvpT/Ruoocn86zHF10QseDYfrjBpDrWVA9Y
h8wouBtVeeTF0eIbDU9Y5K6SeCI1yhHOXbnr/t7Ydp0grG8phVuw22TdyFyQ3e1BZr5lwrBn+yxG
u+8uhSDlfDqFIK4+cMAerPaFTlC+ynWV5SxQiUkRY5QfrYUocIV88shLrGOUJuGbmM5rEh05l1Kp
oUaZBWVgJQiyNvE6PiVxOEOm5fFOPDCeXPmqSwLjVTARlnxgIX5xuRpX9hfPWIy7V+RWbgIcMhVf
ljAwnJLA3nJOQv27ONO8WFAqL/bMLnYlQmaGRtnQHWTKhQoH+xZo3qWIYq8Q/tEmya1erEsaLXtT
WRuJJrmgWQbnX0KdwNguA/f2qhDrQDWOxaNcSorKwipR8OMigTp3pkbe2OC8BhytCXx29Ak+3E8b
XLAnSRCPL+dua9YDUlK79a8yY7/OUxwzCcKDKyhGSjMpa0plmAXPgvpa2Bfr+bVrN3tn1XQI1VZc
/2vTIP9VrMjQ8tTv5sIe76MJzfMyBERxlWHIq4R03WhZOERrlap+/mmGBaMmXTOlFpO5EdIE9QrT
CZveQVQpFOgqyw6L4jyzqzTf+OZnXkx7g8btp0x0UGyf9KtzX1g0cXU1IGCVquBcvuMcga/nYotG
hq8c/LjGY0CTvJr8E7yzXsVhKULGKei9LYOk3Qew53jBqaTo3rfXDUxeROLNZwMC+Jrjx9G8lesW
QU8sldO4FGwsE01BjJbO2f7JHDtGjH/+VdLsJiNFn1pZc/yuSNcugBMwAHsvvpRKDvJimcz2MEKK
F3qWEYvyKHT0tMwunFmp7edCIx9QiR9S5a4aqQJD08KfL7e3slPjhqmuJ2Lz9iueEqqStj3wG6em
5RIFwFGygiwOfdw7+QCnT3QDJQ1nt00nJPbrFXNNs9ZlcvHkIKIcunSO3/M7YakbUIyDKjfnV1bO
ljxsZlJhQ3L5H/1ndeVkJNukH45W+XN66Rk+2xbxPWxvHKBGjKJSZJe+8z0Y//KTVKNOrjz+itJE
l9Q9tS/DymXDXMgFoQp0ig8fryxq8ZXni1eyiBAinlBJVr4sSxpx76Ikh8b6r7VP/LeArG5DNZjY
1M/GdZA5P8d96VAIEitJVDzngBK6lroQOUfdMd4LaKwAwOp9McWvYQy1XC64hQqfEPZip77w44ux
kGrrmQ+caBsk40UjOmH3i51gy4L2OVoT+nu1ThZVRT/zagYl+upkf6RnKklDmbMFRvMr+s29lF5M
wWdFNarvIPRTXdUFPX4tCpqr1oBt8fJPvS85KK/1HHt/fKOmpE8bf1/z9Sd+/h4oSZK7tCijt10d
DpHtdx8mt0782FLaHgZMYSP4Ytk0MrmLfndAn+b6fPvysV7lXyF+W5MHhxmWcuivMG3DPGCShNMF
bqSxujuVV2oZKC9GZu3BgkahxvgrX2NvRvUXr64ezHSgBozFTvmKyJcSyDUaZZvKnj7SdZRxmgNB
o9mz85yHj/tgKE4i76Ys0LK0ncLe388Y27oqmOlxDkTRBF2ftMVsDcw7TJXor6/NJx37oRs6r4Ku
UIkHjMjXAalsGunugE69SQiK6o9NNvhSb8R/0MQUylHgmgH1N254Y/+Aq2WaTe401YnhkpvRx13f
WRrdQuKzBZINi0YDCSOLkvSMfVhj3P5Ns2QaieYk5/OaiWhUV1M5003aUKHvo+ZeTek9rtYIk9wf
QGYbJgLgvGu1t4FHUMmM4l/LQs0HUzKZbETRZJHOaGgBmbP7MHTH3uqY5xcfv8+28ajnet9HoFvC
0dh5RyrmD7NvN5Q557cpb3/0fcFjzaKh8YY+Kj4PnwW+FpBvuO6lu446y1pQOW8np1TowdVmVBMs
O0C89x6IMOLwOrbwbG7coFAV4Sb4xqynPcwlrEgfe6HZ85ZYZpP2mlErEmvveeWzqoPiVz8VnjoW
XqXYK+pPIOlDgO0nppYEG6HoWYYBDhpG7VP9EPx4BkdtWiu5yE+UjSlksc0EHJ6sgS4I5WlewGU6
nIYkBiNVmgs7UkRYX/SgXrpb457ZBMcossZTnYLrIfUV4dojBJcFNx/fea12D34vTVbURsAYJXNs
eP3zCLBiab+KPjB14zFjOpfIBsa0aHeQIgwFmtsvLtbiVQtr9FyB2NX/juS12k+MthRRnYG4NFoP
5ZtlN6k+bO60TWSRygXRJFEBTJazYJpm/nDoaxG4JpXktX0ST80i2ziGOSWL+hozeMh86B7YQfA5
vYWHmXfu6bsK203bVOCGkVcsvh9Uee8LGstv7aChLCMzRXZF+ZSh66v+FCDdyBiFT+qKBhpLONya
HAOeYGFQxvtaM/ME8n8wUasKXOB4HFnqyAvk0D2dKS+liCL93an9eQuNbasHKOYfGBFn4xiYUR5d
HDYktqCb4+kcFifF3Hwchjv5CisFHZvRgdXXAXGPd+bf0qD9slxC3RKHg7TigZAy5ToqhkFQ23MM
rg+4Z4NG9OwnqxMgSGrq8Nb8ECTaq2ty5w0qKS5RMF1hyj1PnQNImBVZqlWQJvz1IT3AJt9vBkPa
q12jQwCNggdpXZBDgtD6VaU5NMATjKdrO/cdpA7myCl7yntFhQSogHeeBvch+XbXuM1RTTc8769d
tZbsgm+TNqRhTelXgilCGhAi8ChYQXQ4ytVYGU8SQy1y/cjc4wyl7r56awVM8hLsddGPBlG4LxNT
PCeI9jGvpuVISu/BslZBQatjrbsXoUsV5OKEoXvAB+mjktcUDIGjYcuYmmJG8I+4
`pragma protect end_protected

