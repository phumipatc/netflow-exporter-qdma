`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
fR2YEb2EqX2Sz+qVm4m0qKD80u5ri/Yw4N3NM0aecG6OASyP4I/6NkqeXXG72dWdZH0s+lP+LJVA
mrIyCernKaRFUV6pk8WG0rJHq6c6UatxVko8IYgXYF87kbqZEXwEUOJua9FFcfqLGJLBqLkEauE5
GhnZX1NCgFjtcReKyHuEyaLrIuUgvcJBULj1KbW29tUCtZsFIYutJCFlXzFFSJoKrL0BNLNxbZ1D
nQ62xZBYuvxUNZcT5swE3hYfkMBJqdLEHut0H1oyCCMq76hhfxsYRdVwq5KEgYeBOh2PX0Ag755z
FZ9bqb2xwwkkzrr1VbfVjrvdGskm7sP+37kr6Q==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
sdYu/0MPlSS3AQZRrL6WYpDNfD0shKIBgfG8HkBYmyzbY+f8i7F745TkFSbjcIS+AWXLd8ZbbbY4
tpFWW/NY/ChgCYgqu4kWmYv3P52rE2oRreEzENscXtrjnV7BQKE2CRbS8D66j+bGpGnFzIcwHQc3
MS2bswboLpcp2l/eo/Fh//872qKwJFe+FbeqmRVooGQrgmD3kJ9vUr9jhDxkvFD8zpoA/QowRcjr
1om5saOddD3IQdd5bdLv83x2WgPQJeSPUi/fJk5PDXbU1SfgPQgjDZsXP1pHY6AtjHu67dksT9Om
zUJWzPCvcqNXALnp/Krh0JmE93f6H8INp4lPEwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
qv90Ktuwm+wJP+8di8rkG/m3Vsxw1O4D33nh35N6kkFSTrqF3zr6hJ/WrRpbMw75G0DuOLqGsD3Z
QpdPHODaAg==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TDMqJ0MzSEXhb2LgxPejz5JHc6mgzOHajdF/Aw4LWiTaiXNr0h5PRsHkJo34VfXg+zzsxMyMQ80x
2d6b+0gwbT8A7cMsEV5+/VtPwwEJbvNGTe2WXaQBQDbqO1grjaD/8RYIm1x0Y9gTBScxRX0d7w8/
xg4uPwaMtnxOUrotHBWkFLYo1IX/bkd5m7osn3mIUBz7+46F2DGtVGp9XfRJwNZHC+tjsKChYfzJ
ox71WcvUjO+yzTkPfNoGAhREf08DyvqBVJ5PUyh2h+WxQXe2rxF4oVePNOFwOjliWo2s6yIcOqb3
1NZEQRVquc3I2bSLOVjVT+un2MNiA7Js+wF1qg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Cw1M2MEVwfMR9ZJHISBfByf59FPflgg/NcXODQLE0kjkxTg+pIp5dFockL/5DP1J80MOz8/IS7/4
QlUtix7xRX+vQPAzEHCj2c3tT6yxbIRLnmCOmPY/nIhamru0S+AfDKOIWyz7ifcqz9648W9ScA/V
y6i5yOJYD4cNHoiYR7QeN0Pjxc5GWAUTeTKj23bUFIOjmryNqcm3zKe5awJPefyjqqnnBbL7tDph
1NPOoK0y8qPWz0iX/kAssKuryeFwn45b+qD2ZHFeJUzUzZdqjXUOClvqMcaTH1wR4KSON981m+ND
ek7zBl2dd1hukaOefFsvv4Y3YkR7hAwcHVOWew==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eh4Ew1q6pon1rpCRD5CbStMBU47QVYEvqyO5nZAb/641o24NesxLkW2NiweY/KaVXoJn8oRl+a3C
fTJjLhvieIhypXeFa5aKr5+5V1tYISkwtpvxLWMkKzEVRgxJTDeYx6ACrhYIlJW1QW7BFaRfTouO
uk1raP7OXG2Fv8PVaP8=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
T5H3zCbVNUbHpwNLwYmSDFEdBf3yPEaixv+PeAdP4lV2/Dra4GjtxJrtITGiCM9hlYzqaWjnmCd3
zt+6pIJ+8iP2cZEng2MZyxe2y83Re4698/CPpjaZ0JrSYIHD1WrwMEZcCehUUP35aJu5nAlFa7zT
sMmP4UNmEgp3o1mB7su5+hpE6t06BaDid3IVaCWVrlcEFm85rPQixQVjSFfmQkfsMVP+knLHH0D+
ix0nhBjbV54UY950XjtPmpwubtBi4SdS2H7PfYTXkZqY/n87YkMhyD6XTxlyNle3U08kfU3L+fuv
924K0b+/S1HKKVgVMX5TAKbmpchD/36UXh9YzQ==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Fw4/YH86wyPeLKJzXUHXlHe6cY1RBYB/nVKETD6YP5206ekYOy+7JqkNRwNJ+SjJxIrYwV4tpvTC
UfCarMoZIOc+r8QX/odVGeB4/4Phwcq6+vPXKWcunV1g8w+UNton7eYWCXWMPCwjpBQyX5umRdlw
ZOY9suCH4QrGAuqmynNOrpQ1mTEIDimNSiKo/ybtB4C8huKZU82ibg8jP7txMSzvEDVjDRn0W+bl
IS2KzfhE6tBPiWF4vrab/FDw/j1SQkI09imEtjUu1mR84r9m1HvviG4HkUK0MvlxOZpL/ORnCR7W
5hPxQZaWawePr2sufBST+3QbmdfsJzrg4IxtjA==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
bepK4fCj0wiD1hmVSTBc0inbrUdHD+9Jyr9snn0SUQUJIc3EzfFJjPe3OokTCQER2SnOv5qpYMJZ
Zk+3YPC5Ev0jXyHf7JhR9xYiunBlCEd1RvaCdZqMH5J2bSAv9gpkDDiRd/GeQdS3VyOIjc46Yw8W
3eiEhzyxcx5gzGYrpow=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MxHuOvUQy+L1zTSxFvDvXN8uN21TKRhFe/NYbD2Vz2HNl3X4W6g3Uj2537X3ltvYtMI4yFHIWuZ4
ZF62EuRMD2EANOX9T5OhCQPsQTpMZDIzD8hvQ8o1kPgugkS1rUlnrHYrSlRAaXDwmXDFoWGOrS3N
lwyk/SqGU4hLPn9Oa5Qho59sSSfyDiIV8dr2pcIzpquddxUbZKVdJavcbMWaK67i1+qAE6tjI3mJ
4fnMqYSqFplOBxF8I9l/tXo+GDhJmPSgTKStEAlgPb26WCV2Cuok8GwMuzkNIb4lbDBuyVxEAFpY
mjwpGbiyWXiK6gtQOmkP9ZPagV1YWzdJWkBZRg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10864)
`pragma protect data_block
kOoN7UpX05Tl+dk08Og89RiEAdupkVzjfgACeGYnpVzLaIMUEbBR1jEtZ4GFOAYcVl3yFsDJNGQv
DOm6F707tKDYJL5je8hxaRtYaY1rkAVfOD0cY4WNOOI4/zDArioW9v/DLRzXltA2VvzapomiMCHF
6vY8yqMZJu9n+aF30hW5SnuB+aDzX3lo55ZDEGvwagOFJPgCLofPG0CkkJzCmHHsAJdd46S44qbR
VWR1/0VK89AlLqLzZ/4gwsvE9B0oPyefEevA2N7uSi0gTeJ6/mb010tCoW9FecIFGjJwr1NFEU++
45Xkkrj0Ot67GBoO3Wd95Btps/W8hxN3iXDeWNrEpK8jbPBKa20ZeMBxT2Qpx/mVC23rGLaFGdhJ
i7CmMMuSXdhSw1ZTNj+r+8JbBVijw+gNtARzheTDpO1cqMhsqrpGo1eaXY4i1MNUKnZDCA8v29BX
PXry7Mc3ed+ENMBWBhi9BXdaoNm3th+5UYBvWzRHksr8rE0/BzX2Iam8mOvj08n8xvOGGT/3rubU
pNAKrzDx9mSNnZ5BQEmohWTaifGColjDt/TU7vlRShqS0UYEFq0O8EexCJbj0MQilr9XretbQyfm
I2n1tKMrf5xnKpqi+czj/y4OrhDHNgKVZpe3DuqCtVgV6/sziWf8TuoahiwNKT+QPEp2jCjRjJgE
RIFRNv2qlB/wTvcOKhXPBTOVJIAsZuNonnSZv9VvaOv4hQvqCVTHxHReE4wa5gMXFnISo9IB1wi8
wOZl2ztQuvkYoE1hBuoyaa5UI8OSn0JoyUQIWZIT+rKKyCiBBOwOi5+Itlwyylg+tiK+IM92LbUT
mVh1ptOOYsJe6V+C8kC+VTQEer5yOiLTrzpYlqYmgtBMvwbbPHr4qqEBApx2BeiEK16XsewYtmM0
gfYgGP3JsH8c99RKjmcn1SFaFH0frWFFfTyUnvOni5hoihrzlj+g8A+ASdR2LS9YkjPPwWJmgOF5
a2x9OIv/i1+OeQSkUATS1M1/TxkiismnKIF3Y8Ap4H4KGlmuKQneNTZfxkWFFkA5gZTs8IGPylEx
XdRxe34hmMA8u7d9Tx0KZx0XhY2GXDe27AR8edK+UBINQQ9VgCKz/R/jXkOHY4j+Uv5+uXibn9hw
M0r0RNS+P3njvUOIWRfp6b7+9WIwigwNDJ1jVbK1hn0Yqqp6mFdB4phu1ubRyOqAVpYzgdTIpjOZ
nM7QpJW8qdwByhwIQEv3z0Q/3zYUPFNi+ad9UohfDXH9IaNve0bl2127SL1jctCIo2myoVNRX8oh
GiJYAgLeeGy3RtICySgclE7bgVtgKE0eYqDzY025CJIMRVSof/gNgtKBN9nqOihE8rS1ga4cFgLH
fCLBx6N9rDuxbKU2/OCPZ3HnfsAepRo7rH+mPqOQ3sePkQfkNVhJIefZMx7UFcgIJN2taVIvjd4y
IhkDNbTFAjyrsC6R/aYaxS9kWyYsD2BsTvmS9jlFPl62B6QMt3Uz5oFj1CoR+RbAMJq03ssmQmtC
FPAhYbq4hxNnQfXbOrUDXljMQTyk/yfWjMXwWr93FcQVnMC7RhEmBxfYwMu/9A6l2o1Ryw4E0ZjU
8k8yLJdZZdiwiKwwLnSKnBWwUdjMOl7oiBpORDeVU8CibK/q9MIml4JnOo0j8OtiHBmemy3AYQOE
qrkD0NjZvL7vOo69VYjZ/kAF2OwzVg91XgVMkxIcnThgCNCM0a0ObCabqpSS6TEwVZVajhkLRW0E
vlDIgNPILV+r8c27TWUhybUsaAM1bs8EigCtbOJ9k7F55AMywyy8qwh8E4HTCf1u25AQvQjudj5B
oZxX1MCq3q1Ja25d4mblmiqGl96z7mczbRS3Y/y3ose6sKuxe5R+n2jM/YSbWY6BMXLpi7Ud1Nb2
Jx2OjFqSyp8xoazjuqkOZPFnRE7x8mbIljHh3F46RJ2XxrP5zth16vWl0I11/aWeCNknJ9jiXR/7
fmJdkNMOOa89hOL5KzrXEMBUL8XjaA53lLHUyTgbG/ZXF9vUArzwHkvfXlQoQ2sOBx07BV5TGUTf
Ydvyjsdl8O+UBgfnn9238kJskGCF706EqWEnCvpGNQtSr8bTPKAT41QOgGtkvslfOpSqPYvmfjs+
Y2R1JAHeR0QYPs3BkE4HMlpEksfNyhe8SjIjjxOKvIOYnvrD78wfk4J+vKxdEqElwQkloFMoZJli
vOO5fJb+kEV8xlfYT7pfz7lWq/CVWiLdKqJRmjIw/pulTtQndcG2Aci14+fCS/eDF3+QeAJSq2qb
GDv8hv5bahWUbm4KdUaypiUxCssdROopgp865Q0nQCc3+GZlln4P9yJ8D+QMzYpmOXA3LaoQcb4X
bVXKhr8ekmI/z6Y/L8cUP3++hLV65mk31nnIcEpRF+vEYhPiBxPVxBNZlVVsxkR8gy+zCzEyd3YZ
yWovuQnH/YMjMHi8LHIVhtQiLwZCnwBpr7vEKFJ1VFMNCNdsjmNwejdNnsCSs/VvrKG0j7/AgSNl
NRHWLMCCQEx+tNHMUQueHE1uZTOr5tw5tZLZZ/rJWwqLOjTQdtAeOfz75rzKQvbWjLm8ded1gdRV
EurXeGHusfqQ1kW4Ls2PWklZUjiBxiqKYKvu6x8piL0+b3QxjXQyq4gSKJjF/DodBxOsNfoZiSbi
TUIGD25QCJ3gOU1C48En+61paEbdHGpwyTyAGeSsaDBbd36sv/jaRcpaOi3MfZv2Ww7KJTfZJ64r
DBfgEf1ukEVd0Y68luWpJ08HHm9jIOwmjTt3XK37wwgTDNOa4UZhPZkij6laKNU3x3uHgD+/LJ57
jaHIZLD++6qgVtvDpzMRogKOXV/VlBEpPxIh6SzPrRYNJbt0jnWsSnK9jZpS8NMznypeW1nl5Avl
DEaYuDp3rxMZQmr/YkoVMX3h0TNr8qOQavzYIcr2VBalMVnHztkR6LKVs5heZ074G7YibEafy90U
vQlzwiXQbyGKusGXELszCkLS4bmoGb/2VT9kNzNuVuDpc2HNCIx7IG/m7+FFCFaL/GbXAHa2p8yJ
fBvrmF5vPe8UWqUa/7HwCqLqhmjwh3pfqA2Eh5wiHgdck5Tgl59/IhS61bqj2Q9jOT17PXF0Sp41
tiDR7JyNhben/CBSOzmVGjowGq8IdOjvja+Lt+Tx0fk4TJt2hnpcouigV2WAboMQZjhX5Lx4RsBF
d/t102hwkf4eRvBS03oWcgiT/GhuLEn9b5WyuYLVKqOdzWXUiSpdcVP7KMwMGqZOjInVA2bMLDSV
/p/xcVtJOQupjKlST3UnH03+jS/zbkPm9cawtABJ7+K/KIen85g1QEXfCXwD9oSxxxtADu8Sb27F
ClgK6knHAaiU+niFzWOcteRev+7ucB8+TtQeJ9pNcCFIdEvjP7NtxjTNW+nICP8rY5osXS1RQXf5
Wq8IHkHbuG8KRXq+Wzkqc/18hOlXS8J6ObgTIxgRiw805JXs+hm9CCJPUdtW6h3hyrpN5pahpmGA
v2iiOBSzMf6EephuUgAeJzxwqO3Ab39TBGTgHMPCtmmNfvk0atsx9lNMiSh4uTtbfbJ3DUGo+Ngh
llaAhzrHywUimXEe6hdLjhnjhOZfhFGBF2SVwCZ6l4p9A6o3J3fwULZYKSaExHbVAhnd3hRjgAMC
mezaxkoPJPOGMuS7KTM58QKQSvpeFkWGv5tBVvyDC36whT3kJarHSq17tDW58u2IRjLORjooD84K
Aly30347mi2LGPhb5mOc1t+5ZPIYNpssLraIMcnKV3MddjhJE+xVd1cyJhVhBcIUr6PrIU7aOCQe
hR7WflFEuuEnX+19yyXZ/ZNU2ndY7JEyo7XpQVcaC2U5W3GIjd0pTyULUnVw/YdE9I0gM6mn4h5Q
nhn6HVyCGLImwUUqlLAe6ZF7Q+D4L//T1FpShzBNQllnyKrbmxwCPuWEQWk91n7SqnfHEpwKNkT5
B0NziBl99ybJHxkWfELBuiC68feOluMGyUadGqsVCq46+j2Afd8ThNsD5PF1XRrw9o4raRqnUQQu
4yC9/pSX87h/qlBqU8BBtcz8sF2OYNYYPU5rL+CJ+QySLBwhrI7Nu1fD9JUL5psZZJ1ncT0B9/Eh
P7dX1ErvpmM1Oy0ITj2NCanZgxbz+l3vHr1bYKUYjwVHD/2woVZcV0ELd8oEb5+rPoRvioT8muwp
hDxz3+7zFOvC26CZpcsKKtNnwTOzd0mF/SGHoodRglX/xy1Gz2bgZ6uPiV0zclGRiH4bSTn0Pxem
x2IjDksAtRFaUXGOWfiXQBWb6BQHHq4kDWwubfUApyy/wlGy4yAyv/vwlb7SJZdM/MCKonRErGtA
eHrmxIirDJhN6sWSuQTuGcz9JYUzDhVFelXjGT/CJn5MeBbLlbhyHJT1jEXMLW7sotVQGygI5YL0
Hiq+D/wM+BqHXQaX/oFM+vFQfGWQAY6v8X95BCbjjyyBslnlUTU1cMf6tOmWwYs3RDTFienvlYEU
DKTAHks6mZL/dpUZtLxixI1oJGaRfik42RhI/3TrKCB8yyYqNDz26yurjT0LkRXGdOG/LcryVQcx
RYSj5bm+qTtH5OoWl3o68uXVME2OkETTD3rfgjDXcWkq8seG2s+FLMPEoRk7seDSlM7ECoykf+hS
gCloJOZr5wzsbGIvqtoLM8QqSpOqGxOe+JmOYGy/V/neo3RLig773iCZxgvGQTGf2fjaVygY3Mlv
FVcbFhlw2BRO9iaIxZ/Cl9vuLMWq6QPKWigjZ7OTdAqtjZP+CvzzRdztvKhoRq0ZEINoZTpPcNRO
2lOiuzU37xI+dlW1zNcpKJoCsuHoAhNiv0+NAUwID24/HTWWREpI5gdxZWhOq/lx3JcOHqLjEJMx
/7wIKxfzXbOg8jK18Ut2mtAF4E3rhaImifVvUSWocEnXQ2p2ELeVOTDVZcFjXZgF0oKUTpAJ2eML
KwWipTiI6dXrjlG2r4XLSQ3I6wZU0SmlEEtxeRsslwdELv9/ZtjoDR3zj8Bi0wPsA7kPDZ41dtAN
H+rV6oXPr5d9aiBNI5DIyWdmzJGsv/aatabHFRafk/z4rfB+L31PcAES+WnbnGTJe4EOGHkVWGgX
czYkmqO4kEMA5pYMUiHSnkqorCEVfG8xnkKD3UEJ13P6AMcROQRMTBnqj40JR9Z9oELDm5bV7ry4
T2UmFyH2z2kIBScwJDJmi3k62B04ti43Yy/p7yHtFssDbrQKtyvt9gtTRcr6fBQDRerB27exuEwp
7D2vcNASIxvDFG/ikeTn/WmVgPNDb0zHVfaRkDggbTjkh1t9YU43eiEvvwo/5qClsqScQHunZ/iF
VxoDlQ+ZtSj/xKOjcat2RI78aGlVGKlLJjogezzhKyeQHLYGtlrSJ4Fo16N6fRK7yDI8KkyYfhlD
ghdm74PNc7YmhYjkogJYTy2f5cBMdetv5v28yv5QGmgLdTbhBipkRmseZTHmWeOzllwK9/7lD9Tl
M3NRRuBDD9B10tB1BYKcDBrQ6nRri1f1QSkSbjV+BVpuN0Bytj7kT3tM9PNxC28KQEkBHPCM07IU
Bla/3fB7FjlbvbFNCZvelw2fMOBjviSI638n/pjz/p8AfGyHHaHFLlRISXbFiR4vGY2YtZXeeUH+
9OZ5yzwerB5kdrFRvJ5qW5npyFv/n8Q0FXFEW/ybDM04ScdNtIjQfwMtJApnil1Unc/ycSjMRWC3
UJp2UIWijuimujBIocOQ44cNs6v7s9egAuQkvNN8b76Cv1AIp2HY9JAb4zk5R4eYbAnNi5gvFi5d
HJMa7yGlqg70PGbaigHrCe7VZc5UM+wO5IL0lZq0oIqZnN4wmjQHKxY2uvlqicFYrp8xNQqFePI0
eAtcXHa8q67P5q71yQ2NauC9pUgAGYbSMNRhDiU2wV3UFc9OiwSuJpQPwsUwtbeIOBDVUgTp1DIG
RovfvyvI89yopq9DQFwbTMO5zhZJcBP4SyKbr+TetvwtjsrHJoj6Yswc1sr0A8OQJgnggrj+6PHf
XqnNn/VmB6ROFdrjuhCvvHiotAtZ/gtsMF/ynOdDj93qrl0odojCiYLuPauAsL/UTZIkbs5kkiyi
Gvpnq+0aI+LN/eS66FNL6jgjh6+FQsJXRCtC4QoPmz1c4O1/8aVCQjw8zSFb+13MzjQ9/VXoHjoU
ZTGXeZ9g6G8hePdNmvDPjO0anR73W3O1yJIgkNuA/DUG+lFgTyep9RabWIzcJGQcmVq4+3FgoZuN
ZvRVQkD4h/u3BBnIHu0ntzElURw9L5YDqYHKyGMrZUo7p/2HZ+YO6zWYY+P60jqQgLMF2/ENwRc9
scOkO7RjTs++ASibxCyAw+MgCv6HslCaJe0vlkRO7dT6ed5M/4m14mzqaP7iTR7ryfD8IsI5kicx
TX479k5zi67dN0p/zlIrlqCvsX6y3sPFdWe3a4cciZixG7ecxePX3wJBrLxWNWX4N4L778I7RhOL
Li7Ac0KM5JsHc+FhSVUvnFDFghcM4ga9UvvSGju64jkD94QyAt4+99n10Ga3wxQUsiyt1+Bu/xkA
wyBmhF5JRgdJR1zTDLOZSAaa+wz3E5GQVb0DGtvyaJiH8XyxB3lQ7vbo3fGshbB/mFAO31LJaWuK
JK9v5oHK7xOVlue5r5pI89FjxjL/RzF8fT316gQOmFRLs2N+wOTU8U9m2vkz3eJOsl5c6IjEramF
2rKWnBNMnUzDsC4C5bRJazpDXWOEdR+FENyvvA44UA6IR6/Et4Z0WwaDmvPu+Fkrw1k2fdFUlpQe
r0kv3V3RRX5pF+kc+xn5jJpSbVPItkqbLxpxLQUq7OLS8ckKbdAd1KflycU6QbLBcTHsPRrdq2zA
adtmaS0Jfnp8zN598pHmHY3lN5lZWnzFXqop5+2RuMN+Hc21vbbuG6edYJCnR4lfa+LG5aBwt7KR
p99xmWzlRJBjk0t3/UAfklZYZToFUHFHKlOa5+9057ad+bnxiE1yzf/y0ULYOL45AD+Yzp/qVQ0J
AhQYEbFTovQJF6I4pwcaM2YEowafZCOnTSwARpqIhmNBGrsrUlTtc7im0JfrnyOfxPckVrGO6a4/
Z2aqiCajc/IyXVPGhkFcRkXRp1YbziZ4YnluRo+3TkmerQg2MF7jNh1mmNAZFau0NRvXd6iWa54i
QUz7cCQpR3dMjk2ShlQPKhFfIPEtlyNzhle3YP8NzY1KPXHKv7+emVPSPjCiK6kfYtCNav2o8YET
hzvjv6MAfFZzalfDVwbWYCaMUwBeEmZUKRNQLroaGUl/W4RGrhOKKmRlcpQxXmboWH2H61tJ7gGR
vpRaraW1ZsEj75uf4xrtRCyOB55ar4OFFlIH4Rg04kd2aQPhRcbZshOI8+c+43trJ2fbRVfPQcYg
yRVAzRGl4gUJ09vrK32whcrAF2BT99R3nh5m1ApCGq0bAsCK/H7Zlw4Gpi8S9kkFVRlG5g377vKo
+/i0Ccd+btipmYItcKiPxlWZ7XvxnKrlAc5WtgRMExuZgth3UQxFIBYasSZ9oNAR6XS6XyYZGcQl
NzJpeKu3CAKxRarQdMP6XMCf9TKmVzyDN0DZyoBlbdrO2C4P1Q4RnipGmgMW7I5D+khLGtw1g7OT
qQuZonEKEulHC4GUjp018tvNKDYJGMLGMiQWaH55jvrQhQ2i3BupwijFPx13GbzdIo7t6EzrVWJk
zeJa82gJNiNb0med8rAUictApcF4POf5kCu5RXeNmiSL8GhWsEqZv/4XD3+4ziTItadQMX+Y0EGp
Ro3fnPB4j5gjAy8IVMvayd4vYbDK2XWaz3jF8xlohAJtoIsGMa3hlOFaGHrul93Xx0r1+ovN4zRv
V+aGy8IoV16bDprZvhcDePyGN9zXaxisAgisW/VUxobSxiHXIWSkYYgb9s4rOsy5XpCPtIyk5hIG
VaN9IWvFC5hi2hmDQ2tDmWvkg7cnk49lc1QoPUMdrUWnfG6/DQzRqU8uTQwpxPpCaVY/UjuG/ods
eELExu1VVJ391jaP1sKRnTwe1rNsfG2epURIN3awW+R3ObzdiE4G33Qxa+xiIbE0be6W0GDibtJy
sKsGkkilI9ACAkafXsjJBX4K9PU6D0b4QTUU6O+Oc434P9Kap2XDxuvM9C5ASPv8O1AuemIGELPb
ozfkdla9YqgYfsyshk7S9QKIOwtGjRj0zpq349m/cItIBYAqDP6RfUIsU4R1XGvdZJ2BOHkz0lDx
lpBASyo0pYAdnRhZ6VKokrMST6NB3HvSMbY1byvpGPnzWtGaS2O4rJdI4vSiWSiULgv1qdqxkWiS
EDaePfuLERfjS56IMeYlzqkfw1shaRkHJ9inLV1Rz/DTlEPWQl/l1fkZU4FFTQ0ynoiGNrQmsST4
QQXfZSiQas/xqlgeAivHMh8ITv2o/uhp5+u8bUvaKu0RueYO2IT9o2AzvG58ip5zqjfedDdlpJiX
C/GxoqFMrsfD02azq7pAq9twxpe205AFCKyAo44htxKJ8RFJJ9YRiET6zSjZz59+Tro8REjzevsV
wA40+Pbq0JJcb7zP4bsG6sVQGB3xp32VgtBNobXiXVZYIM8pMpoyOsuKlse0WoyiRY8Ma6hOaj/m
MTqYxa9UCnwTeOiWwCjQMMmMWjcq1K/CkMp4TF6wSnVNF91n/u32Xjf37q294Du1rKkcAZt7iYII
ks+I469kh90ZJiQeB1iNaeuzoDDC3wZztJZ5BnIpJlhyw7KP+488TZNja0pcXVMndqzUglROgBBd
PlILfHgs8XASeYX5pJKkFKTGQhiN/NbgOrQBoa07obZH1ylGRXH5eVgSOsSTHxNn+PPeSIhboe3M
DA22joPfphrF6mK7VdVOfNZigeZIqvUqNNJy58OixbG1Ps0WQeMr9wm8ZOw/Pkx1RZfvoi+jFrTK
Qpx5apPzAc8gxBI8PFhbhgNSU7AnrrO6acZ1sCisDg02d21O+ZsHxrdBzaXdv4ZQsxZNRgy9vspW
aPVS57k7JHj1nigqnToX6pPdGN3foy3iWRhztTmsTz92k/58nlOCHizdgWTZC8PzqWamcyi45NGD
MxdkIpuctDQsUbTk3uAaisJ//rDVVohUQ0oiVzb4HBWamG6VhNSuhPVIaVAvL1TwVku7+JqDbMLp
eepR12hmDHNIwnFFpO95V1xIt37I7okk529FH1umYdxaJCqOLnJ6T0Yp94IMHyedUQFhjATCzIfY
bzv/tmdZLuvvg5XJb0jVnl/fn8zusAo0eB+faY2J/fKmVA2M1y04u1h07lTaEq2KBt7fS5zbldI4
DF/FqdvPue5k5aHNv7VQC4It0TtXGzAjFaY9KcFEDwGkYCUEzKyR7OhB7H/34kU6RhrUbrkiP0hI
1gTdT7W0TxOCZqdTSt+5736US/2w5ciDYwqbovmwMlgiFTnOzEnp4K0Rh3/YhAoaoeQLRz4Imgon
tsF+JUe3BeTj/5cHB1TphfsWmI1jSvH3Lb1v+pzHToLOpExqV+HYvRc7lJ38oss8L8BvKdDvK04I
levw//6nGK1c0lepXGRCaEgia5mX8nwtaDWoRKpOXaE0Af4V+Trk3wxoFg7YpgkG6goMtpE+SnHY
DZJGjKgW01jIBxJuoBnE4MbaFbjRunZ8UHl1+vJo+zu2k9TlR4vL7kQOSHjd80SjK92kK6qWpVRS
9k7rWkErabpb0ay7xzwaDph9Fw5joxKRRZTUbTKDXnlbNC1JM8KGEkxoXjOYFhihr6c85YBDypLm
EhpLKXwnfT/dMGeHda0vQrfyLgMo14zeYyhWImiqULNrb5wNQXwN1BJ1FfPEsTUO1jtJT1BUVs0K
eVPN6x71anT9UzexsCxVBUB0AWAkEtgsn+oeTBnM/LqhXPeIT/hfo4RBmGaG85aMbgbO9N7eR6t+
a9uVVc4bYXIToJd8KnLgTeltmmVPf43IwYcgKGff5oYsiKDcQjavgePwxJ8ZaZMIqOCG12nRYtul
CWRYXTbOj130Hzj+sQNfV+xfolA6AcqximHWMDk6Gq4blvNTVywE3LREgAHRlwQA6oFjEY2iJtv5
vV5+f0YreNiAR9ps/0ZiQyF6AwvG3NUuKffRKzGRNwOEVDs1vmhM5vEGK+Oh6EvmhpBbDmMuBVYz
kdqEGy44jIjNqEUOx1t3EaK/zmspVRBzeTPgtvuG4oGmkgx8o34W5+jKFGAG+Hz5/dA2p18k5+Kl
iEJtfxFy55eA8Wn6e1Ny7D3dLLMuQtOipmsFsy7qw8bpitmCbD+K+8abqTnmN6mXujDLMBgCx8ZU
7ivwTNpTtlEVM583rYTVTKjxSepp7vFUwEZl+2wAoF0GU444mFlISVES5lNa5n0e1eUufWW3MP1a
yulKYfXUxk9FpBJZCqPJcs/ICXonrgg8v8GBYNXqPh5HwcsPm9TKpPnLfgz6Qfmw8vm+aBEwFFsX
dbHHjjD3a2YduVnkEGiEpbjC59Opk5scROibo/CvC4rWPAA5ihfX3tQXP8aoThN9EUQJi/8Q98U7
g8zHYcZA6xIwPXVznmGChmPBJ/B0zXM9P8Ga9ySB0gM1EB+4XpA62p22lcqixah6+D7jh2l70oMO
Ien+L6c4qPPOj//QAsMwQCYuq7YEgmdwM/UQprbXkQx8Dmft5C8giEUBv1Y6jIaEP0AU8hlKzLfl
PTGbpLXbUC5XGyKnsDvGTlIQMqt90PiqOqpupwureIv3+FhkNF6OrTRW/PK53lbF70ktRMa+u/xn
NLzLxz8epu9xoJIR/aAeD2wFIaBInK8YSIbCm9TMy/KgqzNwrk76gYSd6J03Al/5wS/dna1yNR8b
c7UX9zDzFYYzm6aKF6LfcRQUN9xRAk0XzJjnfHW/TH86IUgDEdBEeSB7thxsZTleoVs9VjOAKtzM
ktk2oHCJ22bIiUDuj3wcvvM8B0n0uV76TmQtbRnVpjcU+jqISss9dBVt7AKDUE0Kgf+ZvWIZv1+u
oMUlqyopbx74ZQUxmqfAUNFAZ3JkjHCHvRn/Mglb/OR2bfGBlqRPVD9gwrvIF/Zef/uSHcyOK4vI
+nW6DdvjqKZeXTsA2nPQCqylZEKtDP86aVPv1h4p4o2oluJv4f7y67kIy1DetcmrFRbxMm7kinx5
6UqcDHGlL1S9rKbRU2PX4og4Mjt9vcD6c0vQe4uMdx+j2vqt7w2COWZZvf56BWjhGRqQ9gsn3Avg
y+UB2ur5/j1p8tDDLp0CPUHGUC1AzZ+EdcExdXRDWuUs92+ccTtPxSjcjM6LXSgMRWp0uPMZ2O4m
O4uTRHrewP8tKaD5nTEgtKJEBzUCo53xA8FFEqcLr6zbg4SdeY1AsPmaNuOJ3JhBeeKiZjoSCiXz
hzD1jGWnf6OiuvVqKUopPxjK2A8hlsiNTMiptFHEbCtZiWRc26cJNgMZjA8e+RsUP0Qmu7C9BQ0T
Dg0JHIkE/kJsyycFdfsk8R1K97GjsVhmAxh1+tpb0XQczeHd/ksVIaBNxtMmpYrZRw7wdQz4X7fy
Qfnko/zYUEtqUTFfETit/YZQMeCt3/LYRRi9vI0HYGAUC1ualSkLcMceH6TMRSMQpEHQYecOiKrw
3yPI9xV+ga4DV/h8v/vRrAnH2n3QAz9bHg1WHpUC8hH890hqFcnbti6PwZwyYVKFC5pvw/TRHFws
rSRt3flNo9mUweT2nkzlzfS8zqfoG/sQCSRdiPjBDqJ4vXd5yrk25YW0r8K99ppnPwLAEBWW/3k2
z5yFeqYr2mx1ZZWvIDLyrDv2llmyWhrxJqXhIKQFHBKg0mRV/36XLbLgkMxGPCtBf2zQO6hrP4I7
cVXwkwhbn8wddTX8iJ99tz09doP68SeH3KgvDMKb3YiKEJhG9qdZcClKgNix38ImRjGkkVoo540R
sjkwL9Sinns6qIUmfqzWylfDThetIzJfv3El0mIrbMA0hcb4eejsPwPvZK24SGG8VFt7n3XieR1a
YOjWk+yU/Ms8fa3KYouwuHzs/+6sQ+5pV0LdVFBcXPWG3qHXw0yHZudw2LKJikxClGy4MOw0XLRd
5jihpGLAKi+S08PZTytd9JWzt9jM7425tTMjVEVznFk71cBnyAEcysdjnQ81avpm07GF938OctND
HnzSfv9VvszNvOH1f76RnWK6zgiM7UmRiswgNwX+DJRWWwbQP+4GkXGp9B6LiUKRg4J60UNskr8o
PZv+HU8S2sCkN/7zOMyeLaMKGsRJhGGsZ71Icjx2irWXXb7DNLUsokU2rGV521CZw5S5HiEKfS6C
mPQfJXhM73skMcfuyjmnUpPcU+QQVreIdkwosV9dweiNrIRfpJKYHSWXzY4w1YwmhO5eb+FqqlJX
A9GleDaclu0snIsq4gx49jB++EmJiCCy6vwdir5Pqag1HPko9iFB7cWI8Z9ki1o/P6+lcwJVz11r
xYDZktOybNbdO7tKqrzf0mgKQ+GRaU90/Kk+0fAWnAG6hUFSoKXtO9iKFByoJMQJojxE9ZijU/BZ
5oAIgbqcDwofQgnRBWvvfBBaVK62Vl/GjlnhO7Y/HDON0xTVLaerpPtDwor8tCKPc7ijpCtOQv02
yGpnS15EYEl5WxEXff8jinTjc+2M6bJnkA8UP20P0GJHRauGtpE3jWkVikuRdjDr9TxgLsPgb2jQ
JWhHDamg7yvooE3DO/Lrx4LwhYMozGQPoaXiVj+3yxKVR2inRje457IOuMLqGJcYzAOXVBSyN8bj
bMDs6ycWpvJ0moO1dk/uqjbp2RCFqI21EcOfZnPIM2l3RgWh5hffwNrVcR+dBSRXWHCszgRezC/N
atNeAqLMvGmRTPjwm/OSC2cPVZa0w9oCDRy4+3zPGxf6MvR8PYSTwnmJc/2bkgWZPv2QEak1bBjw
55qwl9pUDJ1CtauivrGQdl5eZU3E/8H0/2BUWERtbRFmGSabQG6vKHCFToBb9fVUspbDX6QhorKX
gxYMqgRgqdu25+XiH1IgorULdYTCknArhYkfS39IA9w5sAHeOVIkYHErOR/c+4s0rtnVCXFm2Iuy
TjmAA4gBon+vAd4WnXWtHCQJbLVDo309JbFRwGl2W1OFlGeSZs8xCHdHc/UvLyABmkl6OaEeGmDx
fnmAsGXtXZxe45tIVJdk1f6QZV0dV/O3+PKRpZq9/ZAZevQ66aQKAzYEmQCR4Z/gyNdETAgDFqkP
9zggRh9TLvgpG76WmI/NuRsEERVoNYoNL6xwA93GjMqdvCUdM69ivymaMLGd9zbRUclggsNVRWBJ
/GxZz2Xp3VAbIUzavClFuskoR4FZoeyot2kgdqJJ9wIeA2x3/fTH1oMCHEyFL2BT8hR/Iqu3PvRH
D77mM5OELXFItM+JxF5FdEpZFNR0ngGwKjRTnHVkLgSUpX4NWmX3GKP5znyXDFFIip5NSZg+WtPg
Gmd5Fnr2xWMZ6B3fk5yvPjWc2X3tBN7zLRlBbizf90jhH0v6vLm9fgqGA1tLAtapJUosNA9rRgyX
bebCXglPM/LPEX6y/3AxCeU/kQT6FWQ+4u72jIkz3u8rNVMQvIdHRFCCh5nhQp+yBXz69mJq4GVV
4DIqXRRDCDrdLKmEzVne5YPSTFuthEFuZIZcLZ72MoL6VLUw9Nbu3O03Vd79AbFaAq//yILWoHPd
4IU5WsVAI0I/8m/bq3/+oxB5MN73tWfH50FRDcLcdmy1G9z7SjyYf4fecz0mcRmLQzPdd9+OHFE0
6vbqDAiEXYJgPAd9nO5l0VMAqHKWBiLm0BVVOSTSPUcgLDRG4krspaI9+Zzyyx71lqpp6TNopp2+
aQ3eqltkDbrFyW+E1GAzJdmNpO1soSxW27JUHjW80rzr5JzxpIqbN/Xr7p2cPpSIKICe+RVAK2Ml
Gnr+RRfeaFRvbpZ0khSYVC5wp7eoXJGsOhziZ8UziZcgSjKRJXKo4dg9IDH14h3RrvxFwXMP4OH/
6DFcEE5+AuHO4e4r6qKi7ldf9q+HZxBpOyqYg7Q9qAUEiEk9ehYcqPLUD7neiA5SI9YDhRZXc3vM
jy+Mk6RlKu+oGsvi22aaFwLKnC6dEQMoXK3YO6OLPgexnMnLadc0+63G8Sp3P+InXalLPnZAWBYe
u68i6e2P7GyoLRp4yhbUwPkHJizHP5ucze+jM+evlLP9H3UTGZx7QOrTq5OCyv/LAflKSmU1m7gC
ttj8loKnyA8oJZYMCV3OFwlEe0Vi7BiTsCTbYPu5C7HyrUT+CJCbRdfKd5kQCYd73e7h1sQZCDa1
ijYj1MN324zvxc4Va9Ha7aBLQfdzvALIR+LNiPTxs2U6kKDG01t5pU5IFQexSxeFtnn9ZEyuwCD1
GS6tN2qVeNYXUZ4epvzXoQY9sqMmQZf6SYarG/5FAljJDkdXczHGUNKc1NxZRoQYcTPWI8BeAFbe
ImNNpN6gAfXekjVQNgoZpkpikkATUWAbtAoQ43D1XzwlQfaSedcqphbr6D32v/ixt8mKwjtiQ7JT
k1cO1iFC7SLvLtq0V7fkHCsOOwAuhOwiUJIxBuzz9B+72w==
`pragma protect end_protected

