`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WC7Jy/Nc2PtZ5dYxw66SIldMAY3nXVE1YCoF7m0FSWQuACZJhe5CL130z8obnTpkOuh85W+PnkzV
3J3yPm1rupguVeUvmW/MkG61JhC7uNPpTS+ymgvZxp66eiPJxIMkkLlc0oXnZLtm5js5tnF3lXzN
Qw07mS/z3L6UV545Sc2I5zretLGuaJnZogJDfS67kECGhQSIfVUJf/ae+vEomjFAmnQSypKEsA1K
aVeL82Eg7KxVQh1+IaPD46gcPb6tAAlG4GKIBnLrTkuw+/NArVJRAGV17KIywzABNGNF3etTuTwZ
8NYw0LX3Gh+fuBAUrqpDi6vA3CHmVEOYHb4+dw==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
rB7D4h86ntYofJHegkFVgNJplZbT0kYIv7o34Vp8y3wKPkRIsbaFVBvIqQNZbezZ9kRAt4GGJygT
I8axYmSopfGyV+fiegrfSbWYosP3Dc8iDla11UXT8iU1DZsJQhXLHTVUWcgbWSBFbnJ0lffmc143
+cuvuW3Dy2czbPC/BU0GJICGEl3rOl3WCBhZTlKj8fkBZzCL6vjcrtKTFwEaWhz30d7nLAuKpClh
7i2/EtHfCLo6Hbc3ELNQiPqS3/Xd1mXFZdHk7fXM5TRLfjao6+0SU8hVci4LIbYLCb9gbwtXmUFa
cGMm4YL4JxlE7XEjqtIU2wTnktmB2grKac7a0wAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
dqxoid+kbrq/4Y7j5/kqCG3tT+1IpZ2dsjglr2e3NBeprnLJCFbJVO0oIxiMdDpc92CMg+ZQzcU2
xAs6z9UPiw==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nr3lP7QU7DH6n8qQdwp8jmF9NEDkQSdoZRw0bABYxC1XlmN83Fp5cFyFCF8I1tDUXgcKnmRIQiOy
vD+CfKa7AxJVtUbf9+ZyQam0DvMH3v9YgDFJSnTsKSTE+lLZkqYhsL0WG5aEuIZKIl7CZqpDgw5w
vMiO5ISOz4/Dc9sZ3ysQSo3v00cxa6xLW9Y/sR/71ofASpWQTtCDuxqXZYrR+N2ehE08ukAoEBvH
Hpw0iHme13nzLK6Gr5u1FKOqx3Du87Wah5QsmezAsn0/+Zm8xI8P0IP4ZVrh8LbH2op6pTnju5h4
GJfHP6GSr/7cbMPZruZBs4sTOF9rRjGii3rBgg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ik1U+1ZSfXaXWWgVcppxDffsMfNvymal91vdUSLTZsLeW/ItIqC/5MH3Oo7v5JsuBxSOdHhY6lCc
KF3uRQvXhGbugWNJLFbVvAguCuATgTaZ3QxGtY/S+TmJPssMynejthdkKKB11PKo56Pny7J5EQ+9
Y2HmOG1RubgPnxGE6DidvNa3bymwVXFz7+ujYJcefF6nN96LhCFqHtcRojeEU3qghM3mDf79GX4L
MztLUh6XBhGpd+U6+VbxchggI9KAchKOtRyIKONGMn86CXh1QV3lgxQ2TgYJ8/dZHHxr77NVavWk
68yQ5XAW0THUnbWP/VC0I7XJujzx0GAJQtu/hg==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
VKvWZI/9ZRnG+nbBpM9LJt2MPxy9vBKR4bHcW7G2BmqP3Thqv0wvzBVun9A2X8duiczO7Fv1MW/Z
XMK0X1AhM+lrW8OtGtfxvTzOQ5qLzSikr+gi5YPgyC/bWytVjOKuVZUJ9AFoAg0HAvvLodDNI1Qh
zDBXm2YTq6yp1wMQRxg=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LU+Sp/gYiRhSlfxwsg4t6NEsePxZ6fM50XtR/Vx/gl4M1GbyDU3R+9hT3Hd8wS5+CVVSVEXp2ykM
9EauTbqYZnMMLO8CeQhhDUHPAnGVhnKtOIUDAPW7m9FbHl3i7BjWR6JaUJo00Lf/CRB3H7LUWSFA
2jMOfz8BW8fE22aO39XPo01sDPMvFSJJfj603CFHcS9EUvknCCy/kJEJchJwnFNjkrwul+UciptN
+7iBkyI+gL4GwzN0UWLO3m4ulSEe8BTfF136WubqN0Jdu0lprebz7WoZcLpqjl32HHkrxHYDCQ0w
m00Q0Jl1DEz9EleeHY8+O+vkQYz4/vDR13UVZA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
i2Fj/JilaUMDXCAp8eBPUjNvgk1qcrOPZF0yn6wQ2GfNXtBWHx5rSsnaeQ75lQIb4PwhDZ7pS+6e
KduPVrKCHx/W/RaMIm2EVNgAHaEkwdK+V701sP6mSAu2st6YwsAWcm8qk+SeBU00+qqs2jUlaSQB
zPI4iCyQo43mSWXfwuh7pKvAxhl/St8CAQjtC8qnLzIN3V6NIP9kKsh/uO+puq2A7cOE1NDxoRHm
p8BR/U2eyfRf4gOLBcKQnsEiDEzN+XGSFwC/UDb/8EgUFlI/SO5jHr/4NUDJJkDz7txZ6QCOfqx/
qEkKMtzmNTXeIXM8gY7GbfkFz5mpZJAgz4i22A==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SpSjiLzt5JujiaQdBvAG5LjdCeNmCnfNU5tEU3iRq4C4l16V9zJc+Q0Z0sf3CoI7GovxdqCbqcl4
fvrgWKsmPU9uhU0r+Cf6CqsRUZodZ4mLf4HLgdTSxXQ5mOYVkDPFmCeac/W1biBS5UxbAqyn+7oD
a6vwYjpeudIywOt9Dpk=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZvVACLBtgXVqvkWtutoFXAEqaDdd6CPP/AIG7nvbilJV8o/jtc0fmXtSPArTkaECBbyKaaP4OVdl
AGE++TXwRy+dqLxvLVNQZnx/qF8+Z4zXBwM+EcnJ8GggNfsE3UfvHvnU1aHUS36s5x5kociVWe5O
cm+pn2BIeU69DVDNUQ8glMm2mjHZw9PTLeRFjWn0lbHG1BmI5Fnlc1JeU+VoiIdbW8zo8UW3jju0
ODSVuLp6PKvNYFkcA1P1zJdEgHXTMKe6xyb1qaD1Ae4m0aTGT1yqrlGf5byOhzM4IP9XaiWpD22Z
SmOQFe+aftXSOi1NP0Ux6IjTFw7jW8poSS5rmQ==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60368)
`pragma protect data_block
Wjikk+tvOUU93OgrB+/wvzhW7ifAI2vuSEUtPH3zJBA+yygXORwNAn2c0Q7yNLCFxtR/hUXdVntq
zalJKoaA675ET3997R/ZQGD6Ybj98OMSP0AH6Rci8YQ7/IzPsraVIEbR5oAN71zaB0JjTMuWlAJX
S+8JQAcuQ+dO2E/aozaKRzhpUvaksHAKNSmhnDBQbjEt77FNUqXiceu83J/qNpY+JkCGOUMXGMZu
YCb3DIbAlq0mp6y8K2DnOqwfHh0KSRqylcXcGyDz73KTyTeFhN9Kp5S5KUYUfuR94D/OV5dzKWVG
61ISqWaf6vw1GWfULwl8j89okDC5DjXkcLKxZoKOplbxN1ezKsRnVCQXJOnI8e9ZHpbXyrr4ihcI
+i3ctSDZDh2yvBuWSH0o64d0FH8xZWmLKnCyMX1lmvy9hOQME4geIHYL2SDAlimQuG0POl0GylAo
8kbmaAuAik+am/jNNK1+9ymfWWFVxSXo3SBoZFYWf3733j/xW+0vNl7IABT+LKrS+5ZnFM1Lvq3Q
EptZ66wXrUydqOAGJo6Zwjp5UGagRNf+155CIapBzSDLmNa+GMQUcJGVLcS9oyV1k8lxRWbOrJvd
mIdhGGed6Y5lYbMsDI/wmzWrifXVI7siElMYSNbxJeBg1RMqQj2U7iTNMnQA/xZL04sAsQOBdg4f
lWbKA1eWEmw+C/wSQYnmkEeiVYI3srVA9vFMwlQd5u4KemD2eRmgNAfZbI19NYrYDONH6BYVoQwT
Npd5/+1CS/gi0AwdbLD+BxI0B2xzH8RyOvwGTy5PIAtTZOlmSo3+5EUyW0lCwB30uYNeyBaTOsu6
oueXo6zAtxlXVKunQ2RPXAvtlj3vAM7vFm81CXxlwErPQM8+8RA2NkV55vHxtQwyHfqgZ4ogquHk
2f/5gvVON0Ar4R+hAkuU2tj+kVQVxokpxgvHOhc16up44hLwRnRpn68R0LoAm4tlYxgpayCIUF7x
8lgwCDONVQVIi7kh9uKUvx5KEsg0/VSqF4Mivcalq1Hypagwlz9u6JpPXEmk5LVNyrGpHrqTSCnY
M9dQdjIEnpUAHRw/egY2CoHGccLQ0NaJozAkUFKQCn4ws1UV+KFaxIAXKU9KqmODjGRJQlnRs7o0
C0O037+KTzoZWbCFzQ2UdPlSjMh+hcxtcifbAT1RBd1Y7jNu/zEArzy1A2KQcvOdovqKRxReFb5f
outm/JdWp5VsewfVBInpOxCMB8NZwvvVrKU8HfHyBjciTj5PJKJfImpXHDJfq3cevFAuxrFNrju7
m1euAfKjTTO8ooxdVJUwAXO/aVQOYNAmFfq5CKG8GteTaXgZElydvVXxsldiuLD7lPAen+Nif8C3
VGvrXMmqpQnx7+zImG9ORkzBw1gMA9P+5INxH+g528a1jBp2xm6w8aaexyUuhFtX4F4k+0SRR0sI
LzQZHvLt3jc2oFJH4fBzEnWEyFWabZDNjNKEn9TsK3MV+B7aSLHuxCFQvtEeVG26BqQ8jVTPbQnv
mokYzNTeOplQcYWOHbHvny5LoLP27ab3aqLsdgp0AjYTJKa4YiScWw+/VJ6bLmPmZCzy4x46Yujn
hjUd1LZwo4g8sFg9LaaWJp6KLR21qCEptbu3dPwL53rGPgc54991CLJEwq6k8LwlWpwRbL1Kr57z
xWdK+aIA3fIoeYRitkiQnVMjRRTOrtR4ExPzLb2LcrTRfC7jmUM2Ep67RqTF1hDLx1SzonVOAhVT
hc0hwVbxJEjXEzLK1RHefZXJUsqNfY5yHmu4nVTk+XBDavgOLserK3pX4sQQQRbZf9uzKMDa8GOZ
vbgZo+3sjA/QOZxO75mGLIG4bJAKWXKoDWU3g3eQ/k/1Dp6iyRZbI5vCUjhUIuemVitEKj871aav
wf7fqaSoNVeXVzHcyHEa2VaWticWtQLPgK+DotvGed98ulrYefgdkF1lTmWlNIFR0NL4W81bx0mF
JASdbPWacZ5Kw54yQhMBOZXTq0yT2hGhAQVI0uktq7GB/rSo0h9un74sbA8Q8+ErfEhG4reJ4aAB
ELJrvBYPbxie8qOGjKmguZrVx7AzhXQ1wee04dAFwOJHr91PYyq5Qpc9zp1+wLa/xJ0y1xfgh/Vb
ri5De5fhfUldGXyx9a9Amc0XQet7Ck7kgyjTd/ANPkhBF0m/eFd+WLWhg8yJjhVeIW4lsaHe13Bw
Pag3KGdrgJJPEAGHg1K99UgfYK1gAUJpFS2bDIRs6z49Vt4rDUi/5xLikHfds76l3VZexYq/M/h5
8I/KL+4ho2Hu4nN2zI4WtN7iYbPAAtrWzpoAzFWoKRXEHd6INzztdPIoiUdH9BZ3JFU3GRYZMyKf
18TEHtY50AiJGa3KzZhMA2OBQwFsAlYxAESE3pOIkIqNZ/wEPDIsd9KmjxXPF2is7Wd6zqZhQlwu
7AcgHAPL6x1YDmfLDy3R5Yife6OEk+Q6BArwUXHSEk0UEhAaURRTP7QCoYdb1mE3jkB7J9207N0b
b5UrhtEu3GV9YHoN2YUbCmchScwsFCpq4T5lrwb1VRQ2Kd20q2IiVRht2Jib6sLz8QERwHmeE095
BNBDdJF6CFbmu03sHjdENWUEtBJ0XDeSpM2aV1aZvPh7I4RzdEAXw2wtVhlSBm5jnS6Gr0Ou2Hrp
7oBTHPqeYbmMweiMjYavwj/nfveBgv17lqKLIFDEqEAfp4BQQOX7fQRXVoQITfPMia/kOUwAiQeN
088A6v5DEt/WGMSoNJKD3hlyjyB5tYUKUWFAJ9rXS69+dD8oB3yWABdkJDQwPF2IohAUvuXaiUCp
PSOeysVcUF30MSLTGhZ0Q0nUt3bIsnRnKGgN1+QLyvZtiFrHH4MGvnhO2y86wsuHBj7W/WSMnc6V
IExVZg9IDSBeuCLC4LCvQjcNP0JecTjBsfmMnl1annfQsYofE70ySuGpYp/krX65yY2w4ufXdHVf
EqiiRLyQj7XsbRY2yPllnFVwhJnVvTPmlTss8GEmP4ExwcGS9v8W15yI6Zg9Q4wS+C0tyfdtN5vG
XXoo04PQgViM/VHxwBbDz3vvJrXhk5VKqBeRSKjvOLvwRnOA417AahVTFJAqeDtStFOpE0A3rC59
hpZ4FVoIW7tHHqtZnUrlXy42XDcUQ2v75JGKlHVXL64ryP28j1C2a3BehjKFsbiDfyR08cM/FSQj
l91IdSlePwP90rgfRdRcrJnuDIhcNegP7Nw7kuEHcrxq/Xp9eFZRXEmV5KTbphmq1nYfDVdSz87Q
KuOiB+py43akIG2urVi0Vu1+B6dWZbIsdDYBPrSYrfPnhDcAQpVWl/+h4Ie8v2lgWobClU4f4T9Q
6tEyGvm5TPIg3gv+8gzNcDhYXnD7cta2Qpq1+SPIMbKrBpM5VyX4YNSWnqUFkxXcVlGSD64lXsaV
o33AWZD8CSjdTCFd/A4LkcDyY9bCb086G7ScXxhnQwG7eER+NkNwL1tjWECfCv1bCG3DxT6nwQxe
McgnE46dG2XF+Irc4DUi5EgaaqKQVXZG42d4QaaUmyNTe9QdVz/n9shX+/1s0sTZThqIt3FB+nHt
DrjJwhaQazNHLpTIEV0V+bwiEG3K2d9uK7YTj9Ke0nwf5sdjV5wcojrCbGfiZ2zB9bNDtFvWGYCq
Zpyn+e/Os7csB+RIomAsb+goDM8ACEFWI5l8X7vGGvKXXV8TEPhwaGTsG1P4q02i/mkpLoVqclfp
bRS+jaOjEclvkkRPS9gbsn1jnIa25Bl6xT3XOWr/VtKYm7MOnC3d/Lz5ALuQ3DQUE0Iu7cHBayqn
kkeOKbjMh9AGAEYXOPQx9hXyLHGhUKaVPBPOO59e+4Y7hpmt0CItjqL+9MXfPGb35i4aIccz+DfQ
sPlZ5K0xPxQmd/u4zlJj888piaRuhwfMOp5yFCBjPkOjgmgyofPc9pXB8tNf8ZcV+c6CUXK4iGXO
0wKIHw40hMnjk9UwT8Dykpw5JFotUDWsFLfDFQpyF9Zvpne0txahPJLgS5ExFjgrxPPumJKLGj/C
kFPvu4i78y/OOlhlhpUZLKqyQcj0E5L7IQ9VaHEdbi0wvJTtYE4gJyfhrcq05wqKaqrR1FKuXRxm
A8IjQZ9sqWNOnh19v5grpuiyudxVUciQXqrUQixVcshr/7UCrTUA95ePA6r5dOMLrt/L4bTcgs2B
xkNhZxc+RIe22WyktDfAq4+Krn5D6NpTCgkewV6h1uRbetNoVlILXRzB0ew+l/0J/EjiSASAzTmh
HiemQ7YUij1MA33/WcvqKO3J2LZcZ8AJD7CfiUw5en8BH20txQTuxsVq5M4XeB4dc5e++5ByCJ7s
H9IXkh4HkmQMIedBcp+xRJL/7S4ieNWP5cSrftCVlwz2k/dhkx1enbpJXoionOq7p+JSTIlfAPLU
5UUr8YFJ7s+YNFB3cmyB9FzVDQhj8rz2HTJQWb9FEVf0yn/fuP723yaW3bpHuGFZraVx0PIZ4lVY
0GN0iN/FOtn0zliIsLcD7PEW/vT0BOddl/VbZg31r1ZOdoDS9C97DA064zxqtCtd28mYPsqFvLmm
2e6me0gfqAmsgboZ/pbXhlPA/XNGhEtI47Rn1dgmH0f7jbBmQv5NTTzeMjVdexmlODLP1+YChqCl
WT4SuV+Vqnmbt221f8WELSaDIHFTzZ1mo1kb6wVs2sAAfZ2J3M4J70Gglp0Raua7Syr3fcvUPXwv
GAWyr9N4eYBm3rUgIjM69Q44GsF7v13mu/n/Ok/Dh+kUR5O72/7TZtI2wsEKpvRom/6PdA4nbu7g
wRBNbwkhzc1ZQMxSi31kMgFMO2UjXooMe4oG6FQHifS90L+t3jEHoxJ5hfPzacT2AZd5u58uFvu+
SJcMIMsNzy74WTiytvbcp2/g/s9mA5g2gd6RpmE61h9+WH2IkPVzADmS9R7sc5vrWOUBZRuf7dXh
gGAFE2o6BRaWm8m59Pm1TCk52Xci626OSRQKHAFZB7zHl8AsDyNGtCsiBrepLd4EgMK3h5n8jSaV
kSDXkilkxuWRx8me5mhqZiJ26C7TGyK2QgE0zoJr9X0Gen9lhGru2LT9yXHiX5Pid5X3qTYl1cTa
WomdQU0mWyYtuPkIKKKlgb4LywwIr8EEJOa9W//0slOgmEqwkrGgBUG3Lz//fpmrDnJYeIN/Fei4
ckLs76/laRYGZYiyeX/T4IndME2u6L7UHGMj1/MgxoO9w7O3CQ2jakw7Z98qNmHX0RbkAMGDbfkR
z/uZo9G82jIVEKnw6I914qU6aQJUrILj+SW0g+enLE9TyDwu9a0AWQHpyNGrz8f1tDX+sWacsCXH
Wpdd7cDKbGFLcZkvav4bnZ+CWSSsRaQmBRDSg5oKbv2a0ZnfWd+9Cvui9N85XQVQ+zX2JDz5w699
qDGt+DpXIXRevRdaKOTFIDof76L03kaxcBjGD9+S9PuCruA/N/QyT29338aXequqER0NWvSYSqP3
QphTYSIQ+yCbgLRp6BvyhNuJo6R0AFl4/RWfErubqTvCaY/ZvBBj1Hc7r9QKwfB011SMcb0Zb9Cc
W8pxbU2lvG9R9Ykfw1zdyQp+nvSjiBD2nimka5OwzrK10reAGsatFB3WycnAJolsGNmipqARF1vk
ROSQyRV9OumOSE8hmThf6jiw2eGb9Q+YPuk1fBGdGhKcTXhm/1R+qKLgojt3ILHuPXAQKGxGPSbr
HT6zwmfQB4iacP0fSfoxDn8Jghe7chGMzbSqxkkG8Dkwf0K4gfIBOetuKMjbw/2Y3VB4yMvL2DVR
Ek/utppD2piFbp4VLNhxCVmHYhd6LPdGzRmqJudquFnGjSk5K9Us5V3Jzss06DJxnReJ369/pcO+
CUZfLS9CBLhCn8hA9mRKcehf/jJYwojZ1rPqJzu/3hXkcmZlw4Eerc9kNGY/xj1obfPUa5jxLgSR
dyZh0hx6IAkFYdyMttvU0Z+UsOeLteq7ZZ1ILuW8ZviPgChTvPee3h15JBhWhb2mvpStSK5aLpx/
TeYbfmpCzHwn/ZbfY8AUETkc+wTROzqNZEL8Pll488H+27rY0WPmexqXGedm3A9afT6dyR9W8YQR
11lfUj9hfVaCFdAbBhTEdMTgG5sTkGNISWe7i6IwFa+w6n++5IsPhpuqiswZRC/T5xBouMk27K07
G/Mo39I0ZId4j8dMpDQIT7K0+7wVtyCy0tx/L4+F1CAoiV+nGqIjwCRcv7mErpD4DJ5UrjGOHfzM
VvSdBNmJ45Jj2NO6hfdthy7gmNriHTTZ8/gciBapMzwjlRyKvTrqYvY9MNZNDwk9+NyNDF+c+zd3
7szcqbM71sWps4rMqjbTXMEeajx+YywYvZw+JVW3KeNhge1Ltv17v3THFhvy8SFs/yd4P61N7in4
5JMTNnWByzs2q9s+Q5jnhjxHfCw5veGzvL8Td6itLl3ZVQud9bdRwycr4pNv5lGDIL8dlIk0iDDp
y+1pTaazmKXa4QloweKy3SSRb+5XQg9m38IN1FK55N/Bm0ACscG0YiqeBFH2lLNfr+iTBBKAIeeV
SBGmnMkxtHNUd1g2CY5jmQP+SKV4aerIMnrW/Fw1vm1gTdsoXaGv2vYah8BE3aRYzjcHcKnhScaY
c/fAmhXHVNpauVJqqlYhgkIhjrujuDH2/TEDbbHPIvgr+eL/LxZLflTXwAp2RpzXWXJXoO/hNJHC
Z0UDbatPhhleqGvRp9kuadjwUsa6VWYzpP8sWltUfeD3uAy9hRUDm96hT5QUswRCAIGyTdgNJmOR
tazWs+Q2oWSwPOP/mnvpknr5dytCjB9meatNgQMb0xa4pDnwldmpFQ5g8mfHVE0RBRQc2tNb4+mv
voPjZW9jRJtyDX0Icc37nMO/Nni6LQ9KsEGjwdZdFXd4ZbQpz6B+R6Fg9j6C/hQHSrfvvEJqQslL
ZADtlS+52J+r7xLiCH2npMILjdjRbEo+/S1GB5ml7psaVLKGA8tSo2hretpxxlA6BLDEwG+rqIOj
IqP5SpNvzyMeGODRg8bu/pH0IekEBK6NVL9K9Yd6QfpHqCynjmxe+uG2qHHYstvXHsiwuB4o/jpI
C4NplxGn9SF8faz92CVeAciU10RBpFUJcKbKQF/0nb3HaLugicoscjdH/QT8kksEvsZY1cnDjewX
UO2CqWnlQ/YOPOkYAGEOqV5Km0QhNeJi6l5TROh/85r53ManX8RjiSIJuYLwv7FjU7pGbuMPH24v
seH8J4VKKMarcDvm9gK2nF+78+vjBS6S4GtOooXgnbFSGnCm9xjmJlCaiyHE+aW0TfTKu1M2ZJyw
nBRTQ/0HzIr+TsGsFr/1X2c3GVauYw1ppd6LJwtAeUPsjrShCg6B+kSaYhpEYcx8GzgHh26y+r0F
u3iixTWdDTJfRL61gYwyveiwSe2vJnJObK7Hf0EifL2HbCMm4P2IfcdYHEOt0CYkQfrBpiOm7wLm
j/O89yCRACO4zOQzm9Z4F97AYYq4O9y2STMG71kygpSFzWO9T3G73Ps5LhB3CSXqhX5jtv3gFGz1
MfeHDyDMfvXCHwiXUltMw+ZJvpzPjr+SvvHBs5OUQYgn2mq1aiImHjb0oqfHsCcx89e/MXMS7vgr
y9nNtg4E+YE66OiUcirlShaGULgPsGUGF2OJ8vFRB2fjKRtuJmuwaS8RArkMFtPQ2nte2TNwaD+q
OooqCUB2sz1eSD1TLFoU+ZBxRlvXhEulizhsks9WztRzpSW+D5Obbzozl7iJlEnmMH69uu+elYcX
hFhXiyvKt8Bq9DnDy8ddc4WkjVFdVu46IybaVMCZ8L12JA7gnbRAS0DEjc6MTAmT9aZ3T6KYOLNi
YgLk4euFe5O09IViKw3PvYbD0/hgTQ3z+zzp+hbRKCr/1wK8BPKpfqYopLFfbQne35aNISdo8sXT
NiN1TD85Bh/7tLqs0f2wiQ7BhtEnqcxcqHs0FYHdP0Z4u7mJlxBn+88Gohbd5Q8wD6Hd9Fma/xA5
4AKCR8Qov6Y3eKdKYbIgOZ6rohkW7akL5P8KdpLmU89bVUp1VqH/QogmAcrzBNbjrjn8P/QQs8yw
TNpKkcEpGShaHGLV1QsIuBe9kh0fnEwhIRARrwt2ayteCz2NZDwB7FPkXMxm6He1YQY13WbNHfpn
AV85vdkU4QPWitMhx/YrWHmpTErl6QNxXeXFVv4k/BYmjZdGMywP9hfdPLHoJ62oW1fZ9QB1h2bu
uIUSJQM07xvemKl9IjGhRNvDVEiZ9HB1mSwun2Ta8MN1yxAxtnAYPMrPleAe2oMq20zZGi0rWYj3
UhvcIUpBpSv0ES5Ty+mUvE1rSnmFgrCAJW7lBFdKLe8Jwn6QdoclMuoZuoIYwGpuOi8vMkbpvui8
TfuAZQl2lPo40T4JAQl3C6zxm+g9eRMgCtmFDQtGkJJt8mShDSaT0Q4Uv6uwgCi/PiiTzuWlr4NZ
1ZFEKTgbW5Ym9ie5B3JgG6aNVs+GZA9QEZTHfLEtLh9A0I/VaAZqb0wdq2QrWWNZcAUQC+wpyj4G
gg4Xrj+J2u+Ajz9jILdSD9c5LEPfEmR14/nDhEgTlOLWuR14s9gruC+CgL2kxUHHrp5Xahf1HZI3
O02NSaSyL4ujWNz58gc9+2xXrCy9CMZE6E5ktYKESkN9UZoPy3dy85/UCquP0R5gJw824C7kUX/s
A3heb6udw2eDQQzP5NLYvhhRfPs+8BudxvXj6E3p6bfRJ3tJbxx3udXsBlEUdBuG+rbm3vHaba3U
lyUVJbnrg4gD5zqFReGp/OYLsRYcS9rZn6rU7dwBQ4GF63vOjx68TRMlbz/TmDZZ23rX9cxJ10ih
2znPP1NPZGWbQT3euoaM9iEqZzjh4kI4lIE4sJoEST2AYSUofW+IpGGMSXo54pqgSeLqBj81QX86
kcH9nBGT1jjMvbritDOFFMLpVfX3ZigiN5JLoOjMlK/+ZaH4EXbgtrkoQnSeENZxDg4/fluwcfH4
AiIdSPI9ny3O7E5QohsdVC/ZXbiMNC93nHYSSAtynio/pAIst+/Dl9xF/ej+4NhIuM0pBx71XER/
P62zA9kojPiSTNtxirV46Kr3/jxxc0ZpFjxbiUG/8wkCU4/7Q703R1GLijmhmbQAFVGCgbr5ZGue
q2z86r/qdHEXjHxsuNXaH629/5pmDQb4HN3eYI4RLmv4dQFxUQrkvbRcDdm9s5cr+GwrMzoU505D
+3EwGP0FqodT3dWKT25fiE+3viJaCDlqimkwWVZK9/a8t5v/EGTy95kjX2/88Y14oywxGu070+Wz
mmhkQcDhfeacFLq+2121gFWOcXcxnMuXwC0uO9KtMuHH3pXBDbJzGKUJo6XHMjvURilBFYLgCwO8
Fhw3/ms5z/aSuxRnhVawlLlDlsyC9u7JjI80kfw25IM0ouLiASlJoJZmaCAVZ00aGYoTuNfbbf3C
ODK/7XM6emW0y0461/kUW4SUZAXLq/hEqVEez6ZRfBATiXXd1T5YBa3G9yC1lWrauSyLZsi5aYc4
459GOn6OMb+fJWEsUsbbv0Apz0v1cixCiRsRwy+75JwKcAI1pojXuyAYtouKoCuu4d69Ltx+aDoc
qaBjWwjnGXJnYpWNd79rQ0bxA5H3jKVSIl9ER9/8zUzrSBmwtgu3FDEPUlBdf/6r/vK7vcqg2red
UI1PejM3M4yEj29MpLUIdFxXA2w9dmF513gnuNQ74nHq4iVahsIZy+/DDPKPSobY0Y2axmZuDJvW
mRuJ5JvBER+fAPBKeyDLtfznQdE4G5Eq2WfIBveti8iXxQmhvnIEw2famm3taKNjqYCR8k/3SxIr
KMh6+4iybPG9D5XV339fCodlZQ3W8mIw9pL50HqXPXGuF6pm8jX2iRlLG3u119dvHA2Op8TJ90Jy
StQ5cgagyzsWBVPCIZRPD9s8k2l+kZ24zi2+Qv97u/WCINMdOK90X2pG+FOMKV9jDxI1LmOMM/Ok
1sZy7pQUzCFNUn5FauVQBoUv86H6He8lfOKR8+HTPOxbJwL2NlsnvOY2k7ABZ53b2YJlhj3eLic8
0fw1ej82MyyYVo3tRqr1IMY1WHkAats8rpswfHNrvwwh0KhpZqXM9efTS8zdsCLZItkYCdHNC/0e
6TY/e2Tni4XU/hAz6juQxNPhP6EzlqCUiMdeF3VenUCU/3VMFFEuRSL2+vvQcnzNETO6SLy1yZo1
8S029fjCKezxb/rRGnC8PvXYy/PQJ6Jq9Ww+mrJLF1KgfOj1GD0/jGYzcd5X1bX2ec9TTTmmT+FR
y6fLzFM2sT1Tr7TjORO4kFFdQb6wJrcDmT3pcdmVTceOgNszVaKB3m94qaXEdHunO4e5vRcQab/4
tERNs9la1AviLmJAb+6MKCovRwh7fnsw4yn5InNR1JbhOQqeshNjpkHz7Lf+DTFYV0KC5GpyEZRT
hbnAEe2ChiXl1brGEZjvcL3f4g8pkRqOZAlB8SfmxIJTEc8nYcw2tWP7LHI788ZoB5U7jkk1VJoE
EjUYWD6+UUbPXV6riB+0NyFl3lIBHjKoa5U6hWDG9xrhtz+ZX+AP3C8+HN8Ceejj5YkFJcH9Y0Xh
e7ksdZbWSrBiIzzPIMsUKF7bFzKSd/s18RCHOdjofSY8ypBk9FO8wt/lwri2gkjT6BzruTVZ/jSi
e44I719gpz/kPihzuV2Dc9oNIDFUFcvrjFnzQx6iR238uwtGIKDGaj3kandzUhTEa7YdNHK7bJmk
VYAaRCFb7x4rvfQ6cnxj8Vjm0rOSaYipZohqOZ70xYfl9m8pjK2nQLNeh5nJN/69099WzWJvRbl0
AqCyCK91tzJ8nw/0St1flVyZZb5q98cAuomVoMUU/jFPgIiKF3ym9yUd8tK2u8ao6587qCzNVK9T
ECgD+BZoFgUdR0mbv7rZiREGII/QVhR6jDm/Jm6Xs2R7Hy/GVWS28JSlIfXIIELaoXDyhasdctHX
MBPiyv+/Acb512IMp9NoQ8sa7EwEJXahhjU2EU0y+DsX2TmznU9DsXV5olTD67aiccnX8gnnv+3q
iNxnJ8ED/5pJ3WuAn4HXO8GxdFtcQ7xj629NdV73S1hMJ8L9JFDaJqX1E5dae+K3+7hwUOuk2SRq
Tbs+5n3x4tnIDBTvQGD37Y65LSXAL1TXg3hXJxDwhxZVVSM6V2KYD5xhQ3YbEXm9XNlEJT5eEZjW
yWvBzWrQCXIc/Xa8BPo7qKDQaONbXJzK2X9OOWUQuRBeSAsEG3m2SB4viw+BrELQRt+jGEqaVXZh
BT2rwYZQXebNhPENNopvSPbKUXDDADjCuekG28ASNfDjwTP7H0jZNMaTttW3e0g6P9SoWcIUJOaL
U13gncaFTQz+Y8E606l70F8RnLdXrStAspYuHa1tIWVAVbAXYa+K5J6VfJow+5fz5BPovJMEwzWe
PBrjmjU+T3tNLmPmRXpfjIxx96I/JmkpIxTLLqN5U9c9Ca8Sj6NbfHW5tCcP6udIiMAtlfgbNTbj
+hyUNeU3WCYkbE06tWdGTR1IoKZYnVaEgIzavfzzaGSabqK5isZGy/xGdxPK7HRGjPohA/0en94N
5X6MwRvGa3kxLV05rTzT74ofATA+8atLsb9MM46ebF6WozexZg5vcUl6EU/hKMYZpILNwg1BaWXo
dVHlIFbGn1DyjDNa4STNkaPOwVW2QAQJ7J9XS8wEpD8KcGXaTmSexZNAKjrMyio1UmWRIkCmsiM3
S42OxY94Yu7pXCW9AANloMJtfsVPxiW549L3ftIUzq6mvVOaw5HfTs5NdF/+7XeuyNQ1CzcrPTZ7
fNJcgaUFl9o02lQeMsUkD1CAB1cw0f30NqaLwZFm/0/ktPh8awyvE0FIq3M0hVueOFaDUWlkkXCD
fftvREi9NF+RCZlvo/1R2M4bqDbuq/w2TtbJv4CI4v8FeQ4J7YN9G74kBfhwgpkeAS+gSV/pBTSj
cO0vswLO+EB7PkAG1P5C3FTE7cLKM2mTGFASR5hlCqWpUqYmxSenzfp0VAB0xQyxusdRk6+i3YWo
ms7SgDIuYAEftMF+gK3zTw00Yf/gcyHoWWGHJHtt7GpbZGG+ENUs09Vaxixtke7W2d82MEQErGQ7
rNvEM2+Ej/wxZWKJhGXqxj9ieYDhdtS2kFLyYB68fFdSyJIQ5EhSr7kU+nlv2WJ8zMPJzNfmhatt
MlIeKsHzVN+t4igL/tVrxzv93VYlWnred0mN9Q5ks5QSy/JAut2e65SfXp4F07FHrTGgNW0nYvj8
VCuiiUoM3HmUa+xnwH6cATqGcx8lFojpMOcXofYWaYirnzoxRDweg3Chb8XeliRxLggYVgEaPjut
tRDuFFw40wHBn4TCdYjQ/D7y2Q/4yqoj+JoH7D7gWDzbf4CTAAnl83shUtBSi1ohQtNXmJh4vO7p
GVZ9+yWKdJ1TDdWuem7740ImdXkrgdF15+uLBfDtZTMOYamWxrHzWd4vYwUrwE2TJWrKT0kxbhuy
6Zd/t+dE7FGgG8aNfEydyIyKlD3a41Dnsi+NoUVBbRmAMeSBJtUMqDBm99DZ3xf1328puuj3i5D9
EA3vvnjQ28VSezzESdWf+Rkgy2kSpBLIfl5pUz0PVzQVqbIPMPsSoYP2Y4qQ5SHbg+zJoM7JGkzq
D6IsDe3K+hnGQrp/0g2DtjAhW1x2mLsE6T88UlNbXn1dwL5N+6ygdQUfKP8Cp+cp8KlynyAwHuvv
ts0sa5l6EzvlT56nzK5KFVnUYIhsaI0KUebXeW5AYXT4BJpv7gFUi7K07HQaCVuGlVWL11xapFh2
aioitQ60BkZxQSrLarTXCbMEmKiF8ryJ5g10GovFImCQ333naW8NOFmP5MD/pbu+X3/g3QARmaIP
/yGrW226wAfLmYDmcahkwFf9xoRimmyjyhVNFx72OfliT+ZDOVPNYbat19W4Ycrv456ZdbIFlxbN
IeS7Zw8JDzikSxR5NRVIoM3Lx4t0KP7nb2H5nXu+imS7mbQnxz2Dm4i3BSgtx+OTeA/EsqhkZvS+
mMcOGluvI5XGrv6BlwIj4rJVNnGyLPBvfNkx1jEFm1bQ/I/mBKU0IKUWVISqYZO248Uc6ArAaIoU
Tzf9SJeqGprFhTlMZS0yKqri9nPqFjvMnry8VHqD6rkV8KqxO6D3s3X0h8i5HXcMAbWbxZoGzc1y
uOvLqqhmHDMiOiDE/0fL+TGCwZiWhCqP7nkAYo/rceGsoQETXeLZ5ZwE4Zy16OyewshbwlnMJff0
/wsC8O2brF6OGRqz6htVbaLDhBYP+AUOG32MrmkNS0ZyVvKG5d/MtsNqAqPHW+yrdmHZlLGmLdO7
07+LfSk8g83jkVFtwuysRzBlxBc18Y2nXo2XPbahQnNdidj0zKNyfwL1YlSSS0LQ8vVADTU6TDvO
40CNri9WCCl7sA6bdHZfJJUni2osPq3lBwRknaj/Xmqn6C4gGwWMjiVRoV/WmyhobGWAn80tkiSA
i19v4Ez7ZQtGp5Y1+dBWWshzZsrb192RGPGPx8aOEmdIx7X1tBaolBU78tTL0MnViEJ74frIc7EC
EtinFhAVGhkx3mAkj9rQXYKd4iHnmcxCW4YaVcISf/3SHko/McPSKSBbM8pUlpGCf78RiGY9V4FO
du8pVh3KHYkxux3Asddk5TEd2HX9gLAMaR7y7UqK1GRoVQ251/SJ1qPQN7wABa0j323KQf/gCat/
mZbAFPVf1bhlAqZEezoSF8r7wfQ4ZHf09B+AEJcIQuBoOkgtZqsuRfiGiY7fwYF1Hvdps5l18tZc
4oN5NTjlqvw0UgLRAYg+hGFOKHYyiDgCkP0a081v8WysWI9a3k3lHtXzv2SOmWJ0f9OnAXLj16m5
I/7DICLx72f3d0vkIvKzN2qcyO1BrViu22Ndl066BXa6T84LFwFUxIrN/Rt2zLNEu7Qvs3WQOLEk
fjOpW/2vvRtZdWXM0Wk/QdjNjke/dtRGO+7hZjUccxLrnEW5/EmhBPQMcras27Z/56Qv7MvZ0wT6
GNViEC4BZ+t0gIv1lujWpKPMlSMdntVAyDmjLlqLzmFhT7irsPmr/IEVa6YmabH/PwTVEfUg8HuD
f2/KgynDWmIyg70LZuRQKEK+qX7TXn4noQbHNrexygcrmT675WSATqo23qg73M11Lq595CD5zVej
YTqZzQTVob+32kmsztmQQwVpDzRp0owSE4olzX5HZjXEIiHVRNVeEThKI90nMvnA7RIp7SCTk2+x
PsYis2QZptD2v3oxzCfxU2OIqrjR8L1LaMWRyv7dsFEgbJF/5vbQGRZ1Jjm/4llkIT5THICst2F4
q7IU+b7LjnVWhGLT2FOfn9sq21+CXkoHXn+JDvfcInE+A+0DZ3809mifygBmtfzzYHS+I77Yg9n3
rLt7yUtLfUXKTHm6XCf5UxBSy9H/6o5Ln2GVgUnGB+kIm6BO/9kYmc9ln/tTxgHG5+KodKhEzf1g
5LI8Ar8fln1Qe0oDmyznQii3Sn46wPihT9DKVSdFIslylV6gjGW/tEE8TWrRkCaZE0hMD3aagQzQ
0nNzpTXeqZ8Qpbijx6UKpa2tvtxsiBZEw1RK8CWeyOV+vhYyH5hoiFsLJEV8BdyZhml0E6/ji0yZ
294MwgX8jOPw/y1fiPBvPdYgsZlfugAaUsgpX21ETIHvBH16/DMZektmck0cuUyDe4Ecx+IS/yPb
kWUYoRP1rou3Xzagcnjnqex2qer4Fkr4Ny43zLyJ0xWgTXTTyawvstzP0jWSC4l4NfmeVo6/oKzM
NGklaxIiaBIbZz15cj66anCOPiF69jOESs10a75EKnaj/l0wUROIHWIr2dSo8pXveOnslWhwXdSB
OfYvzcscGI3JcOwVkB8IRBT9QKBNkAkwrF7G7HTKBS2R1EcRXkLQez8ZNWKoK8w55nz+ffd5GnHe
Xe19pQNSR+hc5xiq4zsKvwJuLBPt8Idirw5/Ej/4C+zEjJ9JOmF+GFuptCVt52KBriVigpEQEnAn
/rJqZMo+qZM5lu4fNpO0JSTh2boFA+zge6MPuWc3Ix1+B/4JmMA4iI3IzJxPfeix5N0LLQ6htQHo
m48G8i5upF+Out3WXmxTSn2zlbPADGN6wBXyy8hGlO7mWLHiXdCar+kpihH02NiAvva0b34DhlnY
YnZbWbdfd/bQIJPLBdXLIzArQJ6jKOTOa25WHV6HkI52mo1yp6wWQFOhKUrBHgfCUZqI+2IKXd+L
3Sk4nn/XkU2FMIZUtmMVsMbvvuHfcKZjjvI2RI6dbWA771HQJy98Mu1v7+qhUg7bvjmKf5Uu3p1s
zZazpmicnPYZkg5dgpc93sBehzeBsslfKqT1K2T7r7knDxFe1EGvpfxpEHlDhzez1Ydm69za17aM
xHnpaBCK9Hryh3fg/Ipvni6tV99RcNTKGFgUDuKwF1wzILaZF9GCUQv5ftqQMvKdWNXmLyTsAQ9c
BZZ/6aw2G5aFn9EBwqVFMaBgdxdzvfm1JcOVebE52dWNg8zzYu2ysEUkPRI+HiqHWmNQHhxUJOJh
U4BPegRz3Ixvy/HXMAVrsAuY/VlI3enLu5Rq72V8MAvOzez3BXZtg6E+0zkSqKEVlcl5R95+O6SN
bb6pkbs1u0cBAOE4y3Jp/v+VoDv+10KR5EWQifjA2hn+x+oZ0Bgr4IZAcQE5uqSXN8jEjxEz9bcf
YnXfraDD0LfRMc+sQyfonYLg3ZRnOefJQpWcVhAQ9Bm5l+5yCG/lYsUnO55vC1YawDwhzThnlQU/
rYiOfqpOlvndx04tIV51VPbr5EeQNiMMSzwmWRXg2T31JfBcPSJZnKylI7w7eTj6pCWoDCCTRVoI
L3qXBf8d5+Nimh3ZlL1RhBZpEa4DuQIHSZ8Bp0Lml+4r3OCnVk3OvzFq8DiOu3+vvqaYZ4UtNXQw
rHsgdjJgsuJTdr/Zj1F2ZkaaBmVA+6KV0Z5HZI6uOP355enQatVAmhHdNzmGx+1xFvrO56dXnadX
Ker8lNiZ3awL0Bfdk3CDJM+DQRwPa0VwMgFyxNbYku3hJV8g87hWGci0UkTug3wyYox7dX67JJVY
zJweyFxO1O1DKBlXvAaHtNaIawvgHm52UtiYirIWVLuDWJewiIFpzEgoVyz/OO5K0pmH+nZTeDTT
haYYJQBv8AnRZOsr+Fnq+xmpO8Hgd3rbBKab31h1cF7gUJSPaBOYVznWEHEm+HaPlkufjOLPPn9C
VzQ/APCeOQQHJRh/ZV8jKKaYxs7A6iixjdx7dHzdQiY3kwNJiVeuXJZwHa4gy6ouTiqDJedlFuAF
GcM4XLo+UhDzWqSf+/GNu9LFRcrYpZaq5ltdrEeKjVEYLwqvEHUjrmug+a+bJEIi2WcyDnheFOyu
XZ+6epmrYDXp5YyF/mKtWhfhw7GTYF9EIpIvsZJYOFiyuD/zmZY0rqvwZtRguvrLVWdRKdhaIrsK
oKwntcCIjn5TSTtblvgDUwEhG/jWGkUKNw4FdSYLznHFjvVb3CEnRQcbHYTtHyU/wisrIudloeSl
TJ/x/SW4VCTWYqdS+3aIYkwnxw0ixRm8yxtSDpsxlOmX0DReOb7DiDZSC55/LLkiOdk8RiccriFi
cRrpJT8L1z+YBZYYB3kTl2LTeFbZC8/4E9bJaK90wFavH18shTcX6h8jDmiJHwQ7W7iTe9wLQdbG
BkyWaHgYujX1EmhA0Q/8TMRFxWLu28LgXO4lcrPmzkGOdPQZH8hbmGqc9gTeF0uEAx54q0kqKiLe
EYLtK33UzvxIgC9ET/TjeI6SMjGrajUqS/60SxLX4Fdw82onqsKYMCmbrOBuueYiGmX5Kmg1itt7
XTSWFjgu2INE1buavPVkhS5HfgjX/GSBkhMzFwJl5Rp7h1y+UBOA33Lb309+CkfbF+/rrDqyuh1x
CwG9Q+uuXK+ZtQ/y+1nKENFn1mnm+vWh4fNB/mtQu6x+tEO7PW3NVYSdwP05DpZxxZbtn4KNFUrl
R9vUM7cLAYuFPSTQ3Vi4RC3MbZelu74Ui1bZYfQ24g3hdu6vqs5DWS1IDiifm1Hlimu5PqFNs2CD
/3O8A+ql9AIwHc0LV0LtSTabXp796t8ex3BTEi5m2x9xQwWBWE29ZhYGP3GI4k+0E3Or9P3LgHMy
MgmQxnoCVZfAs+hLS2mog+mATfz5TmNgi84/gNi5ybNEnBq1v1xb29jl7vwJoSviQzJNecV4SCbg
MnRsrAwL/MXx8hlBfVnxsegV2eLEjNBjckFmOeAHdb9RRRQxas/qEj2exKDWGZgOtBL9XJU6TYbN
Yy9RMZrblFEIZyHLgVzpMdRGMZew6jipxpLiY1tCrXGYIq4adhiBvPZNQ8fzmtqcGxXJcGZH0YEO
srFDVlDRocVbCzzlOV+ypbUU4SL0ZejJfwFQRTM6ygI9G9v4HIDPN1IvPcl5zpPdJ3IPioLJ2FgC
qGHlJwGw/Pi/ePGTncVUSL8yOvckwAQl+bDxg6LaZrpB1+lNZ6p0t7q1tJCivmaJLISuaSsoHqRf
4Pt/je6H6MMmsaznoRNrruoNSEO1Ts3qxGaPzCeY9iy+jD/dvdXR+3w7iUdMc/J4wgbm9CxTwSPV
GveCKnSY1aHg2foJPilhgJhmkDkIDStlHnXi9UlRrhoCqsFXBYWY9wLK1UhZVji8VZrY8vC3VvaZ
aFd1rZ8pfZOilhJN4VRRf9YlL2eNJ603im4+aXgKr2znRkt1UZv5XwOXYYBxWE4bcpnxQ0NnIKo8
idV833JQMMPSv/Yj268KyGDP+9hXAFeVm5+WlL0OypBt4aPI6JmWHQFKIoN/8FNjZsDCVjg3ife4
Z584CdQEupX5kjth+MfrQloYLq+EVaGp0Rve/UC13goEY2Lq9kD7h+wgdl1bmVACWSEZFdW+5aBV
nQEPa4XUsx/+JapCrcJmqTvwdf24d+j4VI6At/+NYlrmBDfoKhpOfvu5lPwCNglZWW1c4zocucTa
0H62kKnUapeVUdXyV1FElN+50UcUVMJDRvmzjdOGa/DsLcOfFuz9N8D2CUK8NnDaMNtl8a9bf5HV
UvzSpBQTSrk4j8gT/6R8L0uAbQvkf072K54CYGDAsvUUjiVZFHOEngc4OLPnBq1K8ZVBIrwygtZO
SVweUPOMXBwF3QWtOLI1W0KjP7lVL0K6cQ8/OTPKJZuFy4oLmex9xscwFz/WPZofKEFzDV5dBcju
b/ehZDU0BqnigmX+Ubzd86MLjhzrmB6VCq9bzMOAkuTP+6L1MgeuRf/E6FBuk1P/4ar20KIvEtPA
fb00G3C+ahlJys28pk1Q4RX9oxrlpZw0eqLZoL7NV4d/8g8mVGCIPmhPSAjfjvmlSevVjFIRbmtY
4l9pgY0zVjmbGU7wallVpPJylUQvfPuYxnbwqQO4RJeOuNqh3cEg1PKsm0Za1YWDUDRAB24rnlVc
29o8W/XkUAWRqR7wV5lVd9DpEGUu9ANOoLITAeezyzLBXx2m9kOfU/OfGPZXqIucqzlj730ppQoh
+RD0B/ERZSsqXych7RJA/QOTbNhJ2b40jBvJ/nGrRgA5KHUR35UAS4tdVDlYA+Ev7rxUswGTmgiY
CpZsHncWkGpk64Uf4DjPJx/sjWaoPxEvvrgFUk3/v9pw82f94h3KkfxL/uclWkz+DX/WYfk0fvE0
hxwndYK0ikk16Q7WwJy4vUaSmaSddZqRpniNBAXTM6mW1vMuOCy8BH/6/QJfk1Aode7Ca9OxEd19
JBoVkkB+KZzSXIkUqaij2pibLGktzL4rYwIhaj8AMu19DVJkf///0Oh1zL3esuTuy0Yns+iQrduS
dcwRPcxPFmKhmqC1F1zE/IDN1/Lf8Ey/h6mw2u9Rih148ccgea0Z0PgtNfiYpaLjQPuhPTtA42/+
h8MRBGmmFDqM0X0MhGMrQyCKDPXGcX1yMd7fOpq2gYEc8c0fHPONSkj94mGjaGXLzLXoVWbIeD+E
+ZraY4Keatxvuaqq1YJ8x7SgIplQXjqtp9UcqILFOgYDWI8E159rVOWmfPUQaefBkV47uDh7RYTV
/YgqntCt3KWl0VLnTy37LU28dp+IT0avI4i7LVeXvivfreE/GFAYeF3azqvVE8krs6CloDgL6aQl
PvcNloB5+P8mio0dqLIjfDnDRRXFZL7rjFgUWBmA4IbIE0VaXeJxEogSRAV1fG2+WnQsscmSeKMr
kaVrSCVmDOcmbcktjE9VzR0xndjr2Ih+uNNtIgFazPJj2+qtPxbwL633/G/LbtLm769ERY/G6YRa
QW6aeaC1BdMCEsYvf08AnRqxAxA36qkgggmEtwXZauZC79izaOnsw1mGXS+N2EViA32Ae0XJ5y1U
ayHJe+NB+6ziNrJx322MAnk8tjF/dsiq/D464nzgT6g1d9z0es4ZaNK1VAMNzUNMduMkYXXI4Eci
UI2TjzerpFR3oaB6R1VBAklEIvhCt7fU26esjS+CitNRliSPw//8FDcENploA5U8k5oC0y327Zeg
Pj3+yriyBS2+dNd37/0jYUMixG5SDetPrOc5YFtgIRMxITLWieCiUnbJ3LFgINeih5FhuejSRHnP
qhQszUglTt1x47OCYVYJDHKlWo8o+DWnSYvAKhph3ZrFSXxos37nBli5o3HgM3oNOqgzquFlMhtH
SY9pf+FdnI40BhaIbkNbDNekTgEATG4NhU6ieyaYAoCATwK4kMc1k7kpc/UtgckI82PFl+u2/FCN
994dvIZ4KqAS4xusdEwmJvHaIIRjRm0J4mk2XpDi0d76Z/j61KCEuHyVbE6gqKSryYDlm2MX/zRp
qeDB/cNZ/ImJcetD8/oc7mt4+i1VkVrMZSL3U0MM9ChdFt5epoYByWMHJqI8GJum3q2+ekVYFRdE
R37fSpjXKuPae0Fk2VHMu6qy55eIsh0iuw+xZ29skOOVIdkeeqhFBbwiVJmNYEGGGwG/FrmwnFNh
cHwV4OSOuVtlSIjiQTtg/touq61ilyyuHGaXhz5FpImLLQN5fjSEF2BYrI293Zdnkeu2c3nJlp7z
Nnm3PANFk8xlGPCilmEapasxExslETHNZ6yuFz0hKXc2ziVAZpdaGnK1VIDDZ/6lvWBiOZ5yRrf0
OxRKUxkAkkGuNmMsCLM0Hzv3bji0QkVOe94JhnsV+Lo2egD3tQLhYBq0ES0AV64p5tNq/6gPZCrY
0M/17AmDsWSVL8aK6uLTqW8tPMKL6/105L52JnbuYXRqWYG0Vrg3lmRzSCOWA5ahO8hAxmVO6nBF
QBcQT02DbCU4wYeU1yWEWgFU6aevJrPOM2iFryL4/x5sn0bN7RbljqNTaDW0EmtwQSvZNjV0GFCr
34DJTK/V3P9lkY6MiKFJVebgg+bOfDnDdW7kaMCBK8IUK7mTPRnECVl7R14Y+G9LRqlKICDQpsZ+
YWexLgaWN7TusS559T78Quw0Y2UBbcDs9r+tpt4lJSLEbtmaxd7QsPwfPZEX4sMaBOg2EtO3Oed8
Gc41yjkGjk5MQu6sZnUGd/TDpFEhWRgQeZNSKWPtoyACie1ZQ7oIO1Bs/7NLuJ+nyvQWoG3BLoFA
qbbUCJAazW2zI6YjdBLHf/e7+dSe+KaH4Agi/SRECvVBwZr3mumBPAm7nS+IxpI835DWO4GHek1j
yFbXnQTqxYLkvmmUmXv7HUBvzpaVntWxwbwr09PzRo9mKpJmNXnFL9RMlTJcCDt+JTQVMTPfv4wb
1RZyN9ElIEXqq9m5/OnsMFxeA6fwCnLk1yPWhIQ79qXN4Bg5G3WkBuAkmNEfJLQTZfUrgBFCnDsA
wfrDmWpYrnJ6gSz0ebqJ7yE3pDOKF5xwX0AtmDlJxLFCWIHQEQ229PTBpv+KtXYU2csdyTasdoDI
5g3FOtKbPD+E+R7796/J1yPclENczIX3AnbNZeMZjVdRUKQMGuQGNqyRHBQFy+2CIQb7jmCD0EuO
yU/5eiesWK3uPHMu6k6jzJowFvp6k/E19h5ynPT2rN9o2ZfLJi8y9yWN6wtAeovqZL2oeeHMQQXL
zobGrvYbusKb+jGKa2R6rycZ6sL81gERW5Dg4crZyByQCZn5AJlJhCwshl8GA3fSFIcbXFqj8M1d
Nur9iNIoFFk/uMqSjWOPVkpsMNfS2LQmhV2h2BDrrnwwZhzwtOveoZ15y/YgSNC1mW9i8ecPwvy1
uWj/tmqUIDW63lZqOug7HLvOyfjbAz1pZDfkATePgUCEUjl/u8p9PQzewqCeczcn0QYhNt68F6AR
oMH96xBlK86wja8I+aiNYZvaouq6PANiaad/QhJkWJ+cEu6l5w/sRY5kdbv5yjK7OHpslvGveKEx
UCX/BCmd1m+73uQ0eemaRm2i50EPHn/uW4HIcyZF+L4F1THhaa3JbVvm8lhf0aXUrjfCN5w30yJb
S2TKsJHH96IwtP7v3tVVATNbmjNKXyBVgEdFqtuXbhFLfwmDtZAArDDQzngep5XJB5cckAjp0Bjk
U9EYomoxF2QdIGBBroxBhd+Rj8Qay8A1UG3ZqFP97GdI2TmCYrcZazmZdiQqdteIPNOl22hoE2Od
7uiPbPeQeORUHCYBgBFo+UIxkA2lnYD4FdLW6EA/OH8tgdxFPr7Xti6Iqf1oOCqzqYNMJqLvf2qG
k6j5pdIaIBTCQi1ThoDyJK3xl9W3dPrBJ1Q/qG6hxOVCVyWVQeTzj4LF5pT48PFxR5BFiNelxKtp
WM6yzRxAxwVvQgoKl50gXuHMtYxHb8cFkmZ7zQsU5VDle0OfgM2alBRylwprSPmkcvvxRhYFJyI9
vO4x1b+XAaEZbotpIdhvT3gHMbuQroFpvLntx+CXptIEVwmpmsIr+TvZARhHo09k+XvJIrYPFsfz
EZYymUkvnrW5e2Qjj5wD9EnTVS7UUKVUgSyD0gvNqJscDbpd3du0H3yiSS7jBj0uKv4mWaeC9744
xDmJYGQY5+zvw7u4jV9cIS0UKRd62YibHl0iwfL5SqtExlqNVwvaLeIqPCRhU6sZKrPxT3aIlXOL
e90GFxvwvUeteGHtiwdQ68RRf3+cXoLe3la2dyZL5BdxJREteSYbFA1+6CJ0/MupvpFg5piK18Mw
7/UF+/rXzr5YhzjjlHicCssC2K5h5OV1AfTTIS+qWEXvTzkPsSrw7AKPqhqrFyMGuH1e7zm9RRea
tgNF/+C4Ean8laWvxScGpxDZg+BGiIHfPH7+8ufNmYI6w/ITtzBRgZJ7fgYybDZhu3RBwvKgEjcy
z8rtvAKCFsMZI6vgFXOXiWMxJ0WPk14Wi0uvWsP+euapXkI78Le7pSpqwg4z0jPxpYAyx5kSuJDp
q8umELm+422DUV0/LLRYV0ZMOo5qMmtmiCQQrY7pkwSToNb+pucnZuU1Dx3/W3jVGj+eXfLW8d5c
o7AzL8wt8BtRXod86NWzVrDzqnnEgMy0/MDXRWWnEkwDZzi+UoZFXLcSAAT0bAzrdrzpRrJPqQPF
MNvz0kThgXtUKZZqAhYGn6r+eqT5YSl49KEB9cHv6lsU5OU71cED69vK7rw0MRzLu9THn3tT1cMY
tkKVvM8riM2TC0Wr07uwcBg5HiCH+2gBkL81R1uWCVjZDssi7HbZkMGu8KUJyU4AjTx23MFLLjVa
HL1Kq46BQzIJGRhMvD47RpDy+A+FR2rTafO0pChRVqqSGquKvddpOOCma6PXkuYqrxIWlfZybamb
tJsz7xr9Gs0sQGPNqclAYJS9v966eTBp2F5x85bS47guomcP/keSFqxjXNAA6oUiaWDj+jqzbQxV
//irADccc0sAtwZWhv3XtH9eaN1XdKzs2Igw6mMmhW32cVY/haqWbB4qYTMc/ZUF4lVj1jwkds0n
YQWW+5dOU43WeNGFYi8oJgTgKQ1p4JZ0Cr4GvQAsgNeUnCcFdBEc23ce6Hy5YHHk6H+CauQ4n79x
qqe3v1XLpXEXcvV4AT4oBYZuftGD++FqzWYeDYkc3jZ6wrHfzCoX/VSnppNOLjDCuKI90LeOUzzG
tYcMn8ewWb597vfhylfSmADbyLhGZzX8/0MYELwmy2QZ8Jw15QXYORr6tSDueC7yVw+MHwlpJEVZ
bNylv5KHB3h8T15I+DEDUfdgYuaeCiS7qaP9FPIyoEyurqNPiAdaGOxqyCJzujxhZwcULZP3Hsz2
1xhqPOuaZmAqEXOyLgW5SclhtU6Lk306yiAyAwmgiGuERbYQcBoPnvxE7WYjhO/ODgUkaAgEMOKU
wGdwqstUIxIuNwa9+39a58KsHLmQsTOTyy3L9O4TkdhDELna7sWgGeYYxom89pwR33tqShZ+EwUG
SqfHgGg0XBVK864EUZ5BFj18Y2JETlgq5jzzEzBRtXraqfhptvDllIE+NsLjRie5Ks88AV4rF4JG
Go2NXxSYuCkwXhJPPNgUf03JiA8/IvHy28UcC5S7VYwCYbe1v3Vzyut2i5M1mTNguKWP7EwPbDqy
r65Ff2Xd0FHxwihReCUAvBF9h3LA2c8hWv4Yyqsahtl2mLITlEJVNsRUpfIoX8J7RLL597fHYIKG
qQA50xRlXrf0x1LZr7CZExFK/XRNK35beW+WfU7i67XKDW/RXAv6OvVcExAchOEYaNMoYVym/exj
tMOQnwp8U9hDq7dXMvm/2Xbq+9FQbAR50siHIovcxGE5kEUmrHeTXGqUaUdSHfASLDTmAUFTdeW8
+TybBGTSDgBctxfylKFbSmDuJ8NBIjnzi7p/padGQioVkAytma9psSQO+SfXi0IImI5sR9EtiPAs
4bMzjxDdfJl9ikoKk0sGzGvteRq7nVl4VQ5GH8BT2Hh4pIVBnl4py4eatR2N8YUkdyit9UDgdIV5
ghrdgvWqdjbmGYaH7fEW1/H0AKac/P9Xr4dkz3NZVTHogphC0vGIk9jh7ElpZHpn73gwxa0CtXSi
vQxZbwuosiMcTpRRnNtboL+yjEcSDJngNsRyrgNq6rSjj8RI33xzsUcQ2jnQslig41GeJheVD6q3
e+oivsACHDiYG4MZMms0XE04VFnQ8n0qgZGjtEOQ1/9rZnR1Ia6EFcEIua4ZQnhi1oKWHKKWbjDr
PgNYyu2rNsGGdnUIU/cvQ8msZDJNBb3OxqTlS6UXP+W9sXi60yNIhdxubVueVPAnS3YIjFu1Lbv2
wk8Nl3T4Kluce9RoXWUEvv+/kQ34Uur2cvoU/mN1VNnSOzPGjQHgNtFzcHmx6CQ+4L84ogxrcxNH
VRsTpGP+Y4p6XJjeO9CPaOQCFM11UpOq+ikOAERTBFbqPfoV9IntvwWfZCBhw64kvoaVBV6JjovM
E3KAdqu4QQ0znVa/lElFeyqWL1+Ce7yT4/cbj67CzVRrLCx9TQ/JPa6zplBntHAIZFk8TPKQOGWo
RBBve/Adaj2WnSsbNrKadqAXTSsGqDFqpc3CupVChDsJ9TrDdQwXuS+kWY9UmaTk7MBVfLZu/Htl
qEbcFXfdo8zdWImna6oU/uePZaphLiCamag80HqhJdlCK38IKbYrC1fMojnVzHlaXoMnvyxFB7Zq
wFIo55l1a6/T/QUPRyO8Q2h73QF5RWtyod6cvEIv1RE+PsPbN21FulTHfdCEY/Iane+uYlY00XX2
xQXoWinpd7SzMJyzaM7VNddyJRU4GzF6gxdrKYA4cCHCDNZ7viIGTBWo3J3b5pyWYLm8S1FX5B//
oIxuKlJ7pbMYv5yjx2kStcEpklAdul6U/JVy4mmMZd/6LruJ4H1cwKUz/ESU9gOyCQwwq4oJaRNh
PirywIwGHo1SU5WUdXKEp8cfwGTUUn7rOWdEfFdR3h/do+vB6uaBlmkWgzvl86c4e2W2wMajQvSL
N5TIT06X87FC+F4ZMjYM4SwChT5ZJ+cGAd0rGZObZJpU+VoN40vOPRNLVoZrTX3302YahMSxfbOH
eP/kFq5vfBTDju14QFDfvs8DpZEgU6t4ZVQn3YZR/BjZZG+JkZQXrftQZOgCJkM2BjxD3KyxrjxH
auil7zpM4Q149JPHN91GcnL7PK/YmKCVHSeNj+emjNnueW5Rqgy0epP46uiqupiLcm3+ENFWbzhR
IDA89RVTjroFgRuZgriAoFrBMSZeNeSbYY50o7JK3nFNCf/XiPzjZKYg7bPZsgPT1Va1QK6ShatE
9clCJZ0Q6l+EwK45G/EPEgHGeNr2SnKBmyxMo8F5Qei2zoQnmL3Qy37XhKTzXMJhD1TCxKGOF3Qj
9VwBJ4m+0gy37eBXX1iBB+DMBmnACwCsRmgwabbVPdKW6QduEOngy0/Z1e+P3NGiBneKpzVV6AT7
icU0HQ+OcTFInc9Gs9P2ClcQDqE3jX7RcYCsO8LUyNlh6d/6R4jnO5yhFc+fYX23sm/k4fZ5FChZ
8FgGdK8xSZVE6JxqoXEq1e7Zqb1/S34U5OcMjgH4Gb5OuRjkXh0zhI9iiWZEk9phTeMm1JPyaFfT
bgNNByyyX1364+htyk7esu5GGg+zdr1Lpxy59hh6zrIb2LVviljdchEAg5iEzFQqa8Z5+pnH26XQ
I+7sPaOSVpz0QnhkxB3J+o/AuyH9p1FBXCXltybfYoyRQn9PrjL1NsTKtiPTuEEoTboazssPCsDf
dhqKQq82YTLsVBljpr9bRHYzwZ7fs7uBFM9XbOWADL2qwel7KtVSa7nr+WduKnVoHXQGbmisyTn4
O9iDd+/6ONekq2DteP/51t6HUmdDwZ1l5Lpb5zy9J9q6prRNW4aTWSyZ+Qb7LAr+D2OeUzehy2Hi
UwUXsCvRRFdYEhqx78wQScoY/KuNNs56IglonQnwkTu6oZACQZ9OsvhQB5YGrkOdfwnrJWTtvtYF
M2FAQB82i6OzvkfdXvBx5i15DKPXj+QXc7YwhdhsTahbvGpcDDjBq6CZvTI3Z+Pj+S/xC1t2JmFv
81aw46w2VuubBvCOx5tsASTsOEB8rv+OeHiRIVaKiFa2eGA5JxJjfEPUUiuKRTk/+5UoFZuAO7Em
S7IScEtmEADKD1UTDxcxaNySGgovbPhD0XbUl+s/kJYsXnXRg3AZgil/WL+3Ke0cnH0SkVrUomoo
aHTabRZ1y0Sg2knQCn4T9jBKJ/R3LNK6s6W22aq7c+FMhclC/4+Sqx0DReVTLVxvANAd6EvadzRG
qlUVofo/Irf04hbyIShR7cWXtCv7hs0AgMD/ZyAvmSJd+f7MYxGzwq6OXpUpCJCyq4J+TcZUGAs2
Duv4e0kJPugEnNWKFm7S/7y7TASvJ/TpE2uU35WDq+VCDlDqif9DnjbnZUfU6iy++Lz+LGSBHO6B
T0chT2KwHupTOfJ7u9QrLn57ENtFK7aPz/VoY8WtM3esZbi0kQScJ8P3+JL0EVWLmYBaXIe9qD8y
03JxmNHJJb+2pzzKbc5Azn5+C3tGMkvTdObCXNx9/ESdIdIT6rgMzTv5mL42wLlS8LsXvmwPqgoU
Kw3oJDYwnaNtCRAKjQhlwclb7n7zyGPZHfXlC8j/KCc37qLYxYVys8oyl0PVDJ6pFHTX3lvYjFy7
8BrJqhNYD3SsYeVwOFdByhwVAyLfj4yjEGqWdUKEe5nbTwkjb1an2v8EuCskWAV5XQcCVW750gSO
4/ofoFqqM3OWCw5djuTj8xwR9bE1FBA/UNKHqYNO3GCGRY79tAPYoIfvfZw+89mJ3zo5nCvrKOad
mKBtTt1Jb7zz25SigJEY/2NxQl5GvuIAYEOgKvj5TEMvCeqXhoCMSLh1AQmPUi033KfMvvMEHw2A
dk4gUiufHCjVRx1O9NLROI5jmHw9xqlvhM5OnoqUiWnJd/D2pTiOd2mdw8/+V9Z9jv/g1HRzFwtm
XKZPINSKK3B/J1T/75/AgmhxOKE8Rz9k+ra8fREN814E8I8em3ccGNjyUILHwaqwMIsMjsMG1dGi
ifDNM4YzShhDrIiDyenKDIWmeD3cerb+QgEyaQWUOmwZDXncJAWg3VSINDqLBDPPJ0xbfQawtzLH
zfJiOXphiUTex3eORpVJkVinSdg0XEuFnyFLqrB0CgFcIXqvdSB+UARnCCLCIy5vlF9oFYkPML0n
5+GSpXGg5syMEvd4o8LtlfXlxIBexauxRo4UBfm8t3BVTgU3jzE4d0DJqU4NyfLSHp/Sq7zG0Wno
Pv5k3ksWwxUwkP9ScFiI/NMerJ85Gyjs2TJgcz1qVOBJVouM1wbp04ajzDo3mgVMwnPRMZ6f8z5v
F2wNCfQXSBRLC0iSmPNP2ku9KMerPulVpsvjPfyzjCo5qfoJPEs+lnztwOlDlBYSoqKzXfzx26Zv
ayF67chMJp2Vng94P+DRYSZ3cmibWaqrtAzPkiFQXTv1EkvPNDkedpj8BzLS6JjsLwwl/NAtwWLD
CvE+20k/XvX6siQVDcQkCT8w3R8hZ5io8zQ0RViVBO4OEgNxICtWr4bF5i5Cfo6tmif4Nh3+lKbq
KCuO27wq4orAwODpz0RXGcmjm9Q/UE8HervjZehEkHlCO6VyVkzq/2+p9galQKRRX3K/NIQATvIC
oGKiisqS96cefJ+aVC2xVYG3DEddu5KCVxCbOfs0kyTnmHqc9luaLxlD9ZcNhd7yFrEZKJG0opX6
zTtHxfXJYh60CtLBCWdmOfrXYElaPLavKV2ABL7IrKWei/FJ7de829DPJseQ8QMdq2R2ZoJocklB
iFhQhMDMmAeYCDATdjxV7+/WkTWqrHSgQMfFq59yWMIyzAdiyfXWD47494oSr0OvyX0eg0qx6MD/
kFqgu+6m+DCUbik4LX8bMH42zLiYE0m7ki1cfOUJmnof+gT/X5GfD7mm+//8kounEJaPAAIwkD1p
hibmDBLeNdoX2175GuPJA5NfzhIzjhfY4AAvVipwKnTpdhp/c6fUIbWKyZ/4c/70W26FU3Ca4uTi
DU+VWatyRLen7v87f/AqdREj+IDG7/NmvW/euX5/vhXKuignvub6A40Ztg+gCJ0OMBaCMXCqVgdS
JfssmY0PhqHEB/TRWQpWdbwWLZu/d2Sa5n7gSVhismzg3sJCZi5aPRLfhk1nKA4EEiI1YuxISoc0
NLx27wJxysUluhPMW8xmj537phFSnkYK4EFmSfMO3eUMEIL1is9gm9kulmPiLdpd8cSBhywdgVgv
5cmg8LvYw8h6WuL2GZs38ox/IpUsdNqMJ+DxOsNNC8loizsYMnlpvKEZ+ALN0lPrJJqXBn8Y/6ID
NEbWm38trDmqr0jXu9wzJlRPjWTQHsXzBdQW9xy4ZcuZldwL5psAxxV50W7ARwIk/qG55LmuSfgN
xoAvZPEr9m04BZD49fcBdWVooQQVqaaKPBZ0ZNxpsQRdNqNRz4CazEaqDLcmWqXeuSMaNCamOrOD
r/KnZa4c8KXGN7sgY65mpTUDSQGoi83Za3rDzXkUXua3gqsCfED4n53YJTg6fCRitoPbPo03QEZD
PK1JsHa0Ae6aIvxT8gM03yp8B4a9NHUvEdqrIPbeQNr8owtB7kv/YFGgeDY2trGFLE61L9F4qSnh
M7A9u4wkoJ3PCe/yflYIPqkaGE77Fvadc9Mn8gTvr3xRn5Jrzq+pqdOWs9BUIugb5lPwxyU/f2pW
SbI3TctBlipFA7Om8T0TDUkPr9dwNrXFLqGwXHp8O+4xZ1ZrKpR5yXU/PEL8soP1s2oIF9w59qyx
B57sDM14Y2MqzubfFb6wd6UVauwYPvMyE49hPCXxse1o37wqctatuj+sPKqT0+UGN63+fz8rpm+8
WGSauxl4t0Sz43rqabkap5JQSxNAu56LlfzDrEOWFeXdD2diUty9sjGx3753+2TKhpqhqNLSvWqe
ngV6AXiJo0vFtg4nyhtIDsGF6pjO/sIJnjtSp+5RgWQ9wdTXWnlkWvMsp/jzLTRYFtfHlBBXsObR
8mVvC0DPVkTzSbQq4uwj5EpUKiAfy55VT30LG0N3JmWu4Xlp2GeX3yFxY9FR53EezqIyTQ0vYr77
8bRN1C+4eKwn5j0yf7ulDIM9TO9TNrgXDK/c4CMZFa+HTreQZ+6zzlWZ7Y/7zaJrx9UGfRRXqizd
L9Itg2vP4N0qQpDf7b8FfXJrfuXRm5+SaMC+vpkWf8sYsELLBiU4WGbWzxiWloH2J1Ax/Nr3vri0
6w+OOP6TfYjEzy+XT6J4LlE5EVVkC2wQuqCTKMMo2nYgC37aG+/KfkNX8dZh9GE9VxwxHk8tnSel
RF2dyE+Vq4O1uoGBWegXCjop2+BXUcYV1tTqTjWyt1v4ABFzNGERqGKJL4iMnwDatHi3DJSy+p4j
MVKzAFGt0LlcBgFAY7vyldutp4xvD++0D+9cww/X7mSCeCfF/V3yeHdw3xqQObaoNgRG9tmEtg+8
ciMdqFcKhvoc3tb1xDRDHughsISSSS1S7dD2nYZWJdefWLzCmXmm7j7GCJsfLV2KzlrHl6igNZpI
nyxiyIUV1UR++LEgvIV5t/t6F41uGpxTqrGvuPNWJPYaQSFPMp4RP899mCm4wYxRoqj9/EkNwX3+
L+hfVJ2El9ZuL1l8wBBisqWDvnmZPEUP/L9ZYxWjRTDCmCjS9O8gKgJgLoJ3BXUVKsD0nSzOTGP0
rF7/dT8Lli62HhlGU+rudzv57HGOKlWIDztfzM794kUUqThdE0+2jC2tgpF57XCiwNjFK4uwZ1ko
ybuy8VhNAUewK0IiHkmb84AxJDLKdvNay2jjvrv1S9WKfq9sCswYhC0+uuNnHwy2GxmcfOJG/VTz
H+plaMrJpBGx7VQqfFngJeHSk+8FR1YeX7maQLUhfnUdg6L1iFxQeOFW+Jihrn7XY7SCuhnlDyYn
njilBtXk0FHLgPqFOn2GRGhfi3WE4c6w55WlOK6s+HrKvHD665KU1LEP82XB/eEU/VnMoa9rwp2F
h2rpkejt4r2mfeqlJijbuzy6jn9ax10YGq+yh6Psh6I+Q0YQkXfcMapad58+A39uGEkI66r+Sqve
EpjRXJX4XX2A66V5ohYgr4GKvA+Y8JZbu8hMCi1lGBbzCpHz+ELQl6QmRZp/7XZkJZc1QcsW47c7
uCwA17Y7L9b53RjLYXHeSGA928BwQ96MWYtwZRLDfFZIEuoYtmBK2VfMt1xrC+rC0ejSXEcvN0+3
wVfUT209JJIvVmZAu6CQqNZUOLI9rxccrovtJG5IpzaNHKebPMg7eRDV9GLb7xYsdQwG28C50S8O
Q2smDkyVPTmZWXJ6ZmDPjPS00hEAqmaIr2YCGwLqIJTqstQ2TsWCA+5jaLaS2fLTurU0rlAmd2os
2+NUnHnPLLMsJjXGcGrhQbgB7ybQHGiMRXRfHAr3dwOXSKW/+5iKaVD1ZCEW88AjHdf+iLC8Ymq6
a9G1L9k4pGOANOmRGRzquyklzh6A4TGKYsLLZiputQlRl+yxYRT7122o8ooQ8Q2zc8D+ZBoO/dA2
5QPlPwYVk1HxbYJtsZ23ZXlxNx5dHugcbrtfnAp27ITPXtoPJZOiSEolImQk4z6Kbzq6GGTdjvSF
3/2b7zrQWkfAt6zVLKy91gNdP6sIkf19DgxLpdPFernUgfgttypPJFIUeP1XXuDWD15/XQy/kvt5
GOv01IJsgn2crQem4Qy63hV8/M/LT3+kiZkpR2SQoaW0k0c+ieSBIbk7DanxoUPoIOPaP9o0lQr0
/FVi1NwgsRCUNANUjeZJBqHeKl36D4HNNGtuILNlQOvYN9TydtmI+8+iGfy7a2ZnjRFehGmoj+jS
P3hyRzqDzv1kYPpumga5PZM51W9uQR/mSLueBCGG602usqLeQmYvS0/tBlneoBEe0ShEIu6r6L9P
SRFYDOB7Zfpy0cGuKjfjvz3/QgNHFgSWDNjxZV9dyfhPLzEMVIqIqULk7EFxRmlYbNLGDvb0yVm+
Tq8DamEfqx/IK2fUQLD8n89+RB83rRGp+NHmJfZkfVWfR631Je/iBfxKf4WG1k4+O+KSTULAuCSw
4r2l6NVNAK+9zCg13wvruE6sjfRG5CpfX5MxTWW8Znv99CDrum9dmJx1dr9z2Jc4lmplXYmQ7LvW
pWiMIPWKXTwMdHTqSZLMsIAyd3DXf6tXeuknshwS1ozR+ROo8sLVlxhp5R8X/SmaEewWlkpNUS1F
afg52BkIC1V32o5BU3YKvFxjZf1RmjnzyNvvbvA2T6CuVH2f/5ieMo9KcVULuCCUNezOrtGVxuw5
I7kSgvL4j7IDm5rOZ6ZTUUy2YFrfm/ECgKqAFthP5ONEdedpPRInGrGqs3TRE4kOpPa9GCgAErDJ
rbETe6/ca2spCibPIpNc0M7l8Sw1cxAivEnx8JHR6D0905B/iDlf5WGls35X8tXWZ6KExcPRXoQr
T/sK9GdkYV0sidjj7kMW1jKa9uWe4xti4PG3xGS5ySsSB4eDrnxtu/GBCIZaTDvC6qrM65fykA3o
xjhij3YXJoRSIFe/ZmXs7ia3g7NaVwstyDwUbMUsDf5Q3pZNq7pB3ypdBpaJHKAvXbW9KKVwWQ3B
T/U+qBHi7ZpZsjNZLC5iBmF6iLEy0dYA2CqlmpathV5nQ0GPnOoqcYU2WR3sj/+w4+4M7vajeGlF
nLk8hvP/rCfttDbA2pTgRiM4OSvlek8chupwlc3Q55benMhQIP5SlSl5VuMLF8QAcPlodLRRdxr4
N+SJATvnRqIb6AA71VbIRQyvbhqs+Ums+uCnEn+xgoRu1GMnExN7LRHPwZg4L01v2tmt/jv0wCHM
E5x2qFWlxAJBLnqrpz84rhbE02KlOxdsyCqqkTo0h4ALguYUDa1FrYgWcJq5ALrTuzNlAm74tsjW
G/Od3OdHmuDbkRIQ+tKRBNkJ/arUm5mMiF/P1I9tEelpRCC+3Tin3y5CXioHNHAoGURsuikQ1GDn
tkrx2fboLc9zGxvNHnYhqFEKbE/Nx7bwjlz/ggwjGmlKJsgNvq6tyZQ9Pqu8c/2egH/aMdGCMKam
6ZKazaCOEiRnZfd/vPk5RxzgQixQTEytB5BN0oubjcSiAOK217RoNBaGjHkaKofy69V6RB/URbgq
+h1BHzB7taMJQ6UaU4G6EK05kgeb+aLrE7mrHiRigBGb1x+W90jUGLEWqHwNIpbgJMEObjtyKPLr
9Rih0E7XeMj7ka7+aE4iAbThIONU1uw/Wm6W0gtM8J8CaY2ScsXHIBErGZKOd+tEA38AdBCFMz4i
e9A8QomDca1myLRnxnbO0wFNyxndG/OVGaw2WTwrzlaZ756cJp3sZjTt66AleS2catV6VwAB+d5I
Syv9iP32TANguFI4ClmyJi4jjVC8bXxhVrbenHIdIVFbFG2Mv/p3IKK8tejlLKEBMYSXMPXQdoVZ
gQSe9MjDON2fcuqsdSTMKKiB3zDwAX/MFX1ofi0QxjBMEQtgF4TbYZYIMYgFd0ZJeFFzbZc96Be6
jmwrAyiyz3VMnHzQsy6QZhvr0MvjJdDxKgqK3kLzn7FneIrfXhyi5EvD3X9Rs2u641HsSjSm28Mc
nyjUmeU0gRiANNS2pnZf3liFd5z/RypVRcYiWauoaDigN/VPGfjl4v5jYzSJqm5HKWdy79ffG/Gu
9fgtOFtd7iq8i2TxFiPnGzSnG6524Qfl6p4tHTN3NNtDyG6pQ9Bn9i3RYWBn87QFd8oXPEQjUv22
GqLB9ZrNOBzGOOfaRNfHxpZkcWCayl6cd/xSL3trMhWPkREGOKlAEKBqCq9wGDAS/m1qZIq5Sgbk
NeGlKGez1bYNAo7+L2vtlPm3erq7GgTao0L1iOIjad+Tr5A0l7J27UDZQffRl9LCarnx3FfrWAjI
oLTAXa3n9m/nQAtTy+U7fUoNalDeOU7Z5RvHtKi4SsRr/uvS6EufyciFJb15fXMRdOOw2LbbAZvX
Jdr+qMV5ydE7yF/LVPXKVTuiI+fP1Ntm9DSdWvNC4iMYMz+dAbeidiGuRjnEWWWmH3E+ks6arftZ
NpvL6Ohb3FepKIBd6ON1V42U/K6jYZn/BfFCl0YHvev0SlBb9lewcYbSNUn4JXIcZm16BtiS8nTX
CFChS2Is7yWVt3kP8xOVUWvtlzDXYJHGYU0RxspqZYU5MT0qkWXtNS1NCAfz7qpoZRFpE0ZR5ON6
7i2r2cOONOLnXM4nH5kpQ+YTJXAECUK2aqbkQvsU60qfCFsZktvG9SX9Hqxd1+qU7TPwfqiPqbXa
1KpHhu5er6D1MS3/AWuMPJSF/InLf5Tc8O+Foby+N5xGbJU4JfDIqdLHrWCFZzoF2yJ7VsNDZf+H
SxPCvF1dwcQ4aEbfDSISeitiaX2VP0eCgE3wTMWUWa6gGtiBfbTW6XNoQ6XnnlqPRqRdlRhX48sw
0PleNYmAjvZNZeDofh1Kci/PJNsuhfxdOM9W0u7sXzxrVgMOUUdRTSzFXsg1ReolHgJK6J274lgM
1/iTAnlKrzOr5RMb1a7Z+4mDwLt/SroQ/Kkh85aUdno0F3FrgsWt0Ly0fLMcNR/B5gx/2JdRlDOx
15Fm31cvbtUXMWk3GSuO1HymBqfANm/c2YePzW/79hipYFghlt3vyFLBXXiCDjZhNbqNaTVlUcxp
BevMglJDQKhd6nFxLxhKOhKil536u7EzKAE+PzaDjn/peJ7joTxA5X7TyY5/ZcJLqTEJVqPRn6BA
V1u9VkRoP8sE51QdeGcfRRwYDPv8cBJ8lFZPhF+uDbBNnj76ARxmqsFx0l7Chd5RPt8YKat+jMkO
QR1uBPKQ55uJ7fQ3938nOLWNcTs32zk9Fz8+U40zbUdVE2Rz7Sc5zjzYJDmJ8AxEgEIO4acsLk0c
B+KQm6+h2z0d9eAVdddYbr3Zb8UsZXJggZiuSxI1ctkgCsR2UbP1ZAUrmtgNJ8sMEz41m3iVR7+v
bLlAb/Y5VpNf579Uo+SmmrNEKjWuEPUp4mf7cdWQNPpdHZlJdfuW1s7YmSJxQioZwMwyRa/7irZS
YeotypbvHoJe8FtcJZQ1vGpL9vbsRlkyqyp/J8AzPAyjjqQqz0MtqwyosOI4+++BEpFhekXArX0n
2fprhLQLTJ15tiZuTUVh4AzjASXup29mDB7Jv+k9Jb7EcMfpuc/O9J+TzMhM5+ERdW3hJLMgwZPu
HFUShUvUIXW3NFZUnFfFFOXlFdZk/d0VwMJcvbI7xHq3ASsbxiV9P12Ec20QO3psoSomATzzZaTy
P+TyqADMm9HzoI88mdNtgsMwl2tDQiqtinQn+kt2Ilz/TCKU/hUnSr4ZC/ddliKgmi4o/iE5lktQ
ocBUBz1nAYNCF6l8Gabhfutd6yr2kZlwEI/ZHhXg4ooelHKv3cFPE+9+vieqPmCVKedTO3vzJrKh
P5EmnCqjfZOqJWO6BMzkJVMsbAkP30cP2B2F08BjE8FQLW39dXVv/ScrKn5ZBoQGUEkwfj6ag9vA
TBDAlSxeJJoa9kwrjDIQPf6oQ/R0F5B1m13TrVnUh/jDsT4MAfqXwCIdhNO85vN0dv1i/PDHnzr0
c4zyyygj04Rxqi9woDYi6/8jFzESJychsuUCk4bHYIEaBHVQZ3in+vLG5Kw8XKAgg3i2YgdOxnu3
BJYytqMJD+Ve5tK0gIB7VxvGXROQ+UTeU+xpc8/UCzn4zYh/W5Phom3RFaRT/WTt8B95JRHxn0WW
tzqAO5gkpgs6m14An3U3YA7FXWeIW3kLMAL50HCZMo71XHfmaohPZdmI1lRCFZwlCSNHgN0WPPLY
7wufgSCWe5d92kOO8jUJj0+0qHqWW1mO2kJEdhvI1mOiwpWVwTzwjQGAEmja7C8akt6Ux26517Pp
TFBgA2PWakBkY5rjwUmbESiIW/PMWREIjw87yWlRB9+M37NLvuv7d+aqmAGZoX7eFvmLY965nsBR
7lm9C96aylXTlkG4jwWhwJu5RgcZpoBnUMyg1e3X7RPMh/T72icNCRb5BaHXzR80bPbxdLMLn4nq
K4G+/0dpWKn7hPHq+3kURS8F3JF1u2COqEyjH5z2DArFTDA3KFKS7u/a7i+4FmE3clwNksqK7N2B
dehVWPd3g9jFvCHTZz0FXdES+x9b81Idw+0LP2fwVjdOQAf4U68PN3xHM6LdMdbh4/3AXK51a1Zm
gtMz0E3R7z0QspR/qt4YGEgrhZ3gocKFAVXNIcFufi5g2og6Fi9gitYoDZW8C+FIet/cGDJAMeTS
DRf20TVbmicJsJejLDZZFZnqBjGrMXzF4NQh6UctyBZAuJwFc2jctzM8SmEK7hKkfrMPgDJQ0+xl
k6BPhXxRFCgjUPTU5XDHCFZhZNmoc3IbCDXm85NE6OO19Qq+r37ug3/WSMHYmeNbIKjTgp8cGvGi
1/bYnl41X2rhq2SzE8rMhQoNT/pHonjXq3jogbZAlDOWTxlK2E4DgPCcpgK5NDlsXDLg/AcTTZIA
oGirtEg+YTXx3iN9ENCFCQqVKwxPGuuQBuRukTK3iD8VaFc86DygNQFQ0y0OmaqA44XlhsQDu2ur
oL4WDFU1yqgF7WYdfWddzIBL10ygLAcLFG2eKSlgU2bjiZYEKkVxNEE0/xC/LPUQcYwCRI95qQjW
pC5Gvy9TF8nAthKZpdfKBylZveJindbeJDd7d1H0/1HevdB93+khSM8IycOJ1NCjUQgJ/90PLhJh
Gp7pUm+oaZ3MOiRMZ7qFXCz0D12eyOZ+Zm2AFl/n88dHspx1U6yhR3fhytgom5lLCV5dN4XQWUmI
5nGLJcKjYMt1RPEnVRa0Z/CbJ9tluO2bTf7wjrISMx8JMbpqXzSfe3ehd80u+dRHw0imFe7J5JyL
lFey1l0dsAfp3gRmzuRelnjR9RVmbWmQU08EfRUF1Y86gPsagWgIssSqhIU5PXNZpvUNE8keQdqn
pwqVM1R90ZOZtzNqvZ+vhyISsgmiCmJw9ZPBVKJHhj5SpMQGD5KuLBDTQ6MPFyHnQZT/qX1klwOM
JFJAdSe/pMkkW6d4y0Irg+iJhYgCnTBGDWddhOcokCslykpnnjaZKIvyzNpz/NJ+sUf0RrMbTCEa
3HzsdOtsffaLHloIQXgX1t4r/uSbJsuNCg5cJ7x/j9UZejFdE0p/kJll3hU+DcVGOASWuHeGN6JS
JPmRvu7Z1XWVI55kIkca32E2JlbuvYh1D54wTPTYUzRfXck9L83pfariJOXRUvDsHfQDlE95LX+N
qXT1XJ1gza5HE5yaEZlypRHbLtIfN2BUmRcp4gZlzheEqciZxV/XNM7UHBJzQ3hG+cxuXvup5nmV
wkN2hQe4vyIrPd8HkdbPh3fTFb2OJZdY1f3tLPa2wCWTVT1VMyBmmFV0Gbl1Zb937Q1G+y+motyR
/YWxJreoYMvafbm6xoLpTibhf5r6DvI5G+m0hDmxzJE7nSq/bU/3XyX47WdHJizzFUmtmAdxecRN
303+aEVMlc0Z/HzONI7YNIqx9ghy2PieLJAP93UEBT3HYynL0mb2uPzhaz6jVG2PiQS0PBBV68vL
IP6RTuE/xAobmFenB0T5ceM6w6CzUYfvZ7fgHzezcMLF0f/eZFcTK/cV8ldAZcU5ZTyReseH9Jgi
3yJhLtmHowCqoCJrSgdpDtAtL/8SpW4r7GHxl2ifdu8PRXFGwEN8TFN8+k/1VJtP4GssuWjSjjmE
zhXRA8zDpQKyOhQrz0x+Mle+FWt/oN7fuH6n/5An2rzGLXJAIS+ERT72AeEbnVZxZ1HPksFNDKyY
DZyYkg6IOd4R95FFzP3k3Kh0zH65PZ97k1nmhzC8lxtQgpxx1T0hmlFOw+hQxBo3L+KdNX7JKcd3
6/0sVndetjvtjWZ8spG4oBzsVZ50lRS4kzgHVHzllSE7yCEHrpMDS1r/bCdEe+ucYlA5KwKfKaTb
Vt+rXSOE9RmvfbOsvq1TQXfJn7VACQHdoqsxeygRwyoev95VFzx9f3hatjbvUw1FVgZs9hXKWQuY
poGV+AUXLKH5JjzziyJvQnbhByx5wHU4+akOzDBWqcQfemxV1Jv/oOgx+KC02IEFz9qdjel1+tKf
voogTvvDV4vOB6UilpAkq+n3iTQTjM6ekb6C9GERl5CdNQROv8ZbjWK9nKaQ8497qO1t5s5VfIxC
VBPmZv4JYZbiYUQv9Em1qFOGnRE9bQaQVx742FhkIND3iWU5l8eH4aM9qc0OvuK/tfVeZsr1S3OE
T88WEWoj4oR86vWdMrgGwY3nL/uagkkel4/Yq12ppJLPBdqVnaYzWcdjRJym2L/NJ+2XSJJUIyo7
5lXGGH6cRwRihhxkYQzblG/Ob1SVLC2MgdkrgUCN/E8yOqTqBtjIX/DHEbIPrGodg2lnFjlcRPL7
14KVli597C7UJuzs0MRVPZFtW/Tow/YCy70+waQnXsmuMCa+VqYaLZc4B4GvDHDUnG/CuKNprSQA
6x0TmrQXh+EMlXdxq0836AzdGKQpYIoo8hLAI1Z+VQKY2+Epltff0aEG7l6xJZgoY3KqX+hUuG+q
6nkZfiYw42XLkiUHLy5w1g2A1Zf/1xW4Fno1Y+ay1jGh8vDOYgj/fF+HRv6oTS22XX/JNbymWF9O
PoCl12jgXgO+gy8c3isAypgfXfyZ3qS53pUmuW4/wnTOwUOrOv4OtJ6DZX8Vxy5U035rz8dp+/Jz
rH7bPEBgrpmE1SeGRj7iPZX9GJJw5AM4NjxlmHgnfRhbyXJZkbRbAqahbA36qb0OJXWw9YAghUQX
NnGgJy8sWDq76jaH/TRxY+d34rXQyzSgWAPxNWgqC1KSWXs7MeFQz16f9GAtQFwsO5F37R19z7vr
/+ayPn/Sy7Z9igs+VaLQzxmHyKxlhTEOhgcHWTep0fY5ElsP6C+2X17tllYGOZVFCuTB2BWwtnSu
jxwXtSKwsKuHqNSFkS8RUwwzuBZXGQHirFCqLAfRFkYosVvujCOwy1Vqitw/jAWJXi3jlgGVkpDj
ZkOcf200Xchfervzkq6n2tW/lfcGk+1MSa2Rw7B3E6YEW4JFAdJzhie/wnapfSwXnyUkWB1LSKsd
Ce7dKK9fnAtxpJE0Nk0nYeX/PbboJ63hwW/4pFkAPMe9qkCs5wCbbwJzOos9AA/3GW++DwyLffcu
wpx5ap5Ntzc6N0G2kwDYIMlgHfwW+k3EAArPhFClmBVrM7RU1o7nfYy6LRe2LEXZkpj+efnHgvIe
8w6W6I5HNVI0B31FO1dz5YBcEP2/id1Dpkt9y4Flb8DqpybkESrw/XtZavphDDXnRrIjpm7zYgX2
0yRZ+X2eEhj2k1u916saHfwx9cYzldOCn243T6W529G0pGJGHjT8gApX/+mAC0kvoNvwlnvbi/Q8
GaUHH+dMDY8lPcrySisv6Ea51UWtZjHTRp5HKbDiWzUCalb9pFBmzFHEC6Ks2hUC1I2Podhb8ney
pImNcZOlu4XqljyqglV4vd0Cx/AL/ePaHE5Zz9GMmqdR4gXVx75seKRnwx4mzajExkpCSRcHRba7
cb7ntUNee9PeII17yTb0PKAomZ8tGQd4kvzJuMDag0bK2rrpyWiQkoI6CIjmZItuDsuWgG1lcQ0f
qLyHoLMzSxl01Gjlr24gVsSS5JP30/J5ZRDMYvwtgU+L3bpGxvYl5pAqHqBtLKU3J1IivqUEnGDE
um1N3JGUC1+4bcU2KPf+LDbgSIN2di1ra6jl/dPVCAGVddrza3hVd+pxOw5cOPA7juuVDLW8jVhe
l0HrCncVQO8/HlhMKLfdqHuGL/TPNtJFJyZU3JQFzbJ75iwtx0+pgX9X7gU2ERLCfR6tBtoM48Iu
ZvMOrJ5PuHSqjD9W9rt8fPGBhpVvdsWzMahqvIOz0SJaV6xUyU2RGhzC8g3AeAUPwSnH0eOofPgT
MUqi6ljXQu1+9gEm7bW5Fuwh+/71L8r9LkzHDcq6VAL47TqChH1JTNyFUdnxZX8YCSUVfuv4BZmF
7edCAQLY22vA5Ak0HYMy/hgOH9+c2fJvGrEyDHlokoQfCpGxNM3pIW6lsQWsjez+n1+8KHmcZ1Y/
x8LVIIWmF041XPBSRKPlnO3m8h2kD0Ze4o5Ji1NUJG0eyPgCrFHoro7OoXSXI0KpgPIQCNWt19Al
WIipeTaiGJbV/uRxHD/CvU5tWP+AG6Sg+IVc4lJ0Nd4ayIF+Nl3rurTOzT/I6MG+uOvBMcYyfpdo
bslgt4XQcR91O4D2VVLEGTRR0GZNG9HeemRKHP+ZK47xsX9jiwzfrV6zYg8+SbbdotkX1xCSnyDy
Op6DkuzKgMo+sJXv02P//0i8UDvXMVsBbRrynZQG9C5BFKyYM5mYQqCebJhrRrJtDddLf6F4ZdS4
k+lJZcUYupnMwbxRB5drHDmWDMDNxB27bt92L4hAbqQ7F3izBlCV4ippoD+U1xhQzy1LfrqJaY37
CbC4zGmlPn+aZCrFvEmtvDwgZ02iH+SxFHCS8/6AaV27kfi1AcMwWnChUpra/WhtA+bwf141z7gj
LLjPfV30BaSne1kpyXPTfmSV6H6r7VCLVHoOOc3jYFPnQ2iIk2ZXWIs1Z0Rx82bmlCLIGHl+Yvxu
c3Wh5uJLxhcjlyHC3C+IV7bGVMn3eVXBDsAenwHkrK9fc+2Z6W8ULfg1tgTNPVd5NjXAiw83jywz
Zh/Eb9sFplxGKiP88R1AwdbohDxtH/I1p8pSrLIy2aHFoqxldf7rjKMdPxye0qXH4AH0qaO1nUce
xY/Y34RZlhvKdvGqpAouoZ+fvakOIa2tmn/SJo/2Mps0nr5JeCMS9BgL8vmtxGQPDpA7RZhIE8nB
mMiaBJZjCGr027wTwVyHI87yfy4k2KNsgNgnuOYjP3rtnIwoGOG59MEvncYTAylsFbl4Qme2WGT5
YZuv5MogL4ROc6eghqTtFoABFCAsOYoyasSmts90D2HB5kK77W6+VwCRbVDrvr4iMvzf27gaK5ck
TYAVxN1zq9UY1xCOdN52uMB4M6nqWTwoFUW1KkczWYAI5EbwTWFqVBoeUdHehya0dOk/YUxp9xrZ
+WAIygnJZFOTNb1IfYpzJNlJHqyuYbzbLRi812VOYYxgmoTaOKuQ+gXLlJlVIIihzd1coX6XdZBn
Pf3/Ac+3LRUfd2n8FXItPkGOtJedjBE5QGAi7eI/GVLu6NdXGRu8mvQBfqLWd8zIgZ52OJhgddmd
vNLMEdis2dgVAANU4fuZuQYcaNB2HFQqUXvCiQrCkJnVW48HNOU4H++YvTQcj9rO+6cL1dFSRJhS
tDX2JpLMIh1MWmv0G+SlD1eAkpxdazThBS82LSBWk2CVcD0dJggNqxdEjryMgUV4xc2GRVGoIfxX
S0h4Tc6b440L297pCoe6/lG+/hVDnJ4hS9AS+WibQ7nKnGqo8Xqp2Lziup6s0OZXXQBhP4sDwdEC
XrdkwbYQQWMBEJB4Y6R58dWwMe4RysRjbVJlpeIAOqE0JQY4Rf9zYBY678TFdFEwEkTorMmHDpM+
hgBEetwoOvPmvAmbPLrsaeyR8+YPAmJ1ZiIzQ7WnwMXwXpZrBUbfTuXRWJ/IxoJwt5JYJI9kTfye
KKlunJ8JlGzSw64QlVBvm3T1+Ha7sYOylrPJ66akFFMM3l+TdQyQvIsD/EuU/b0N5Xgu9yELqkHs
/nO2nGwI59fC/K3RdPoYkttdiCRUFZqomOmxTUW8iDoGo5IEx1p7pQOs5Xj2jVbMPBvy168haRNq
I/fKSq65xDltx9/GoEdZt+Iet9e4O7J8dc2EoH7dvsvzCgPen0+Cd/e2dP3hJ4QZbkDwWUTZt1lg
3iWLCB9DTqBEFwp6/xmMshUMYd4yF0A435G1suXAwuMcxDM0Cufo011d0lC+wWt4Mb43Fsdvfxcy
bucOogIGdjpKuecP6mNdI1ZI0ID+MV+t98FyCd5J2zK6IatM0wLWiyML+YQEUvMP3j+lu+r+ME4W
mK09fu0+mCyLb9XcujVYq+WLZa+lA2aQRSNA2vZPtvBOFQ8vT308WhwvbO6O4d/LXJ7WWSJ2/kdy
D5jyoIXsU4ZRcai7TMc6sWJL0XYRo5dpYwMDA7rmoMnx//oTluEsMNK8d/AzF5BWNLyrWM++3MW4
24G293nEU2u21KN3b+uFNMgPKVoMWRGkb1o3I9mo5CjNMEkAZ4WC0ELNBV2VWdzWntjNirf9P4D5
J/3R9K6X1puklyu1x6mSvVuABR7zJvgEoLnKkQuyGO0PDFwcX1ppMFFULOQRyvOICTYsIuY2AT0L
+9/bgliiGCVvl1sGEOhBpCK/XxHZpRp3ZFOiksM1LeMnhwgp7zHXQirrcOK7kkToKv/c++Jhxc/J
c83FI6Qkj/Vub6VGImmkSKCymIaM5D/uk7t7jEAR6oUAe3n8l+1g+wlD7jr/ujxEVpSJdoODFfJb
Oclpo0h4z+WPu4lOMTCnVcDtuECNTCZ09z17LQMb6XjxwpWodl4poY6V+IHP6bgUedYzbFnJtp4D
PESvhGvPDf7FmPqKBLBYScI22qfYxNoQ5C8QduW7qG+qY8PrhhGnYvsp3Rq3MI1Ux5Y+xvGZ4BZY
q6OLC2XKxltr3t8EpCp0v9/mNvwF76o1EmTyhuVgrPOPf3Hkm438oEk1+amL4WMypovZvrfzRTSN
WSzyj6jKN6uV+iwrlVXz9nw4SSX4+ZGnulr8Q/f5+C5aY+qbFx75bFtbnQsL9Dc/HvfG2SKDWEj+
d4fEISvfHZwvPUf832ADcGjgdzLMaCBA1CJnxFXw1iqALvQaI95J0rkI63XeCKfSxyFOBRMWIb4k
VK1q59LHx8uoccq96BIph+JJm5OvXEjPaO4Qq232CmEk9bXjF/d9ki1oZT+7vNZLkqMHtUWf2Yu8
TYiQF7SYB8Dm+fhiCATgY9OB5+EnLyyzbvmikV8h7fqilutjuKUJJKYfw6OsY5fuqXv3rBr3v9GU
6JlAZUGzrkPuzPCbLM0kizRhCWoAkzVL+xCo+C90Zv+fuTpsIdPU7HdsbxGeX1WKyxAuFPEiYCnd
q0CQJL8WiZWdo2z6Jm0noebj8XOKn6lcZ7ZIW1UKso+dnUu+ISGgCjS2St01PuWW8+8lo1FK0nDA
bdtMoe94NORIqLlfYAmUBMBL3nKzCgfxfq+vAAxHfpTc0hiXa7W7UYoRMVnm9Gfs4y0aGFPRsyd9
jZSnBEJxkOjt3W+Geau+cA+vbxcUl5nCnN3DJbI80WEcEFS6L6b9x+nnGTrR+jNgmTvWLeFh9a1B
KyB3mYWxUGefnbmxjBEJkQD9u26VFtU3JEY1mhlzj8vJDjzpFvdIb4ExNYPghgCouteSa8rR6Qh2
mKWu5ejssRGqb/bMXDa+MIjUWH2BvjQslhCNJ4341CHRb6MaR1KdOOn3w1yYsJa3g4H8V3IE8mSc
eEEehiakxxEvVDXcHC04Bqtpfdwze7dCZ7qkbitQ+/fKN6OtXT9O9zVtM30VHsoaTK0W5FIteAst
6Z9CmUiIFlmiY1+k81NI6pm5feo6BaR9o1B4ghOnIQ4VCGR+b/MMdQzF7mrSK9NuguGR40y4Juql
Cx6xC6ixpRv+ZysGUrJC2iL+RCCES8QqseSehFDY8hcH+RYdW/oahRmn6yIuMgRyNwgBXOAdWfn8
621STBjbSZtrKNlFnzL8Ju+Rszdz9AKkWwcHRA5iBK3/6uz8RBmswRaIPAHcUiHmdtTbRjK2Gfjg
I7t5Gf3HDuKhJAyptc4l7bmk+pKHlJQ913f1Z1sDwB5EfLF8vhxyuHy67oLmvKS1eng/S9sAExxt
r4PT2bkvSPI2Q/dB53Oa+jSc89ovpc5YhihLCOz/w1AHzC2vvfwxhX6qjmfUPZeDVdxOSFRw29YR
aThmXcka0VHZgIX6DFXX3nQ7iYxMQ3ngkwhhE+2kVGxjLY5dXgt5mrGWs97V2P3ZmT1pGrDxMAS1
Qjaz05+u5iGplSMO81SS0RGhVox79VRKwNmLOYGJRJ+2nckUk1DrDw0b98UnN82W/hT2ZHM7TvSc
svIfD5YuQwIOSA0G7g1wY/KaT9M4QM1MVey+UJsOPNZZKCFurdI5iIqfuGUaGizBxO1h/elBuUvf
LTyTJUX96IJ7C2xgcAEhDfu+wVR9Dx9buclUBf8jBHIzFo9WZppUSHYSjyOv82NVCJHBKGOMC8Pb
nXM2E1QEyW6l8rw9flTAn5jhnDy5lKvStTxsMP29luw4YEFEtfzvKanjnSfdchICkowRzXdxnm+9
DLJ1nWB/3/5+oO1EUzGip5lILZNA53B/byL59/m7V2xIR5CX01rg0+GL4+vyKgUcT6BOnPho7pdR
sS426mM/K3dwOlqQaxfgsZFydvbBC5GIrQuWT58c7sPZ+HmSIv1UiZ6oEel5qHCwiPWurgfpPqXe
wEig7TaEjbbCGkuZOaFFznPpz3wsbqkRW/fxRz9LanI5FvUsVANIh130hql6HsJPITK3oZLnmh4w
WbGjK2tm+TZbry2YjaoZj5r34p9BcfO8LcUXhgpgXbC/rrEFh8jR4Paijr4ipvHartKnPANs9KXt
hRLPkIYm3okfucci+SgwucpMrqzmJvLSE1/0z+HeHFjO6j55P6wFcVUAAM/Y5nK13RDLBG6o7Rma
KzaKNnPwXeuYk2WZ700CfeFwFArKQi3/XEOJ89czEFE9i1kCHG+drFyES82oiOqdH68HRMuEBPH6
N1tyQW+KaawoArxpcy2uZYAyTWnwIJe4uZ1h7kryTULi0NxtajPOpo+xnLZvJN0OxSQhuJPpXZsh
4O2Y2iRCFY9bWT0QV7qJfnT/JaRwa4GSHOkxg83gZO5RmLA2u2/VHkqD1TcDwMKauiBTmg3a6B38
MCyyq+vgp3m7Z+RDKaAyFR3PKh58NMZdxrLoHb0XTtf7FYzgx56ZTnJvd0nCoIMJYLfp6wEWvvK8
TH1pmQ2AZy/tSNKxnElOZSOSBZ6J3hfumsbl8+36FaUY9+ZgaAok/niL7iU1sanKqdZtIKm9Vpo8
vuox4AuoSvtSRn+sd0dlex/3QlRox43+ZguWws3UIuf4dSwmedqA1FBPJtH8QRdzfYTwL7q/dQvB
OQdTWk94rMgKuiPQD2G0SvAZW0UASjWix8ieEZaukuOkikrK4wFa1fP8tBJ71kMuJrYdBaaX5P9o
z2WejpLUyWsFp6q+6DLfc72fGgIQvtHElvp62D1lp/nfIsFDOhPTXImlhbriuJ2XfkzI3PoU7Cjj
/2V8Dh16icLnLccmlPmPkP52YZcPR5/LDh5pjFlvFBHvZk93iThFnZU8laCUlhA4XULH1PhkFPNz
la4qyKvi69FEibwvItJjtIRoFuOvn39JfgX7LT4ZW2iEg7LvQqKcd78NkUH4d8ctedK8RZRr1mkV
aFZdeoANe1iKgt0Y9pdc+Iu8QzYKWbTN4PGm0GjEzCWBpG+ylvpo0CJGNJCNDHYy2ztvmI7qt9wC
1XONIT1ym4pNQQyk6IOuszSNQn17uggWMqHHB0bmoK9eOZOS+1WoIItKAuNqG/HWVgADwUwB28Zi
00ddDdGr+Ltz7CfDbD1xO1YPtez/02qevFUhBv4X6keDXGaY1Cp5DNpSycWdBdMgOZSuzoXu9oer
lIhAAoHVDqtOY3cTU7EJ4uyWvhKU0qV+M7iDt+BE5w0xLslbozN8+iEEVMLtzpL8LOmQvQ13uSOl
ENisx5qPv5WHlRiF2YM1ap6v+kBMs6xKM6oWcKGHzqq7qltz7Zbn41W6rhA0bnW1qk0vpu2tbFd9
c1NDD296zEfAt8FTAuR+All/AYQD6hljH+v6RB4e6kK4ufO06TqAJiafhrqWZ1B9a2HdLIk1ihvC
HenPCMXqdC5tZ49/aGURqpf4Z5nVxGnL0QUDCxdKZ7YtaAXVvqalkLHuJhmuzTHJOC0kREE9TSBo
je7O6o2Rqe0PX7VgABdhRoeSzrt79uepfWQcwRKsbZS6RL6d8NYb44jACoPAZ7qjj751wQcjozEN
eF34M1UpvRfvlWpByrfzMACLYtFSae34rhClClCLCcbks4+fAIWP8d2vXMgq5tlQVYZ+U9iOzDWX
WlrLQH2vvnNwPzg7mbySfQHwmM+cLmJRqPUl3Q0jhPdiW+sLVajHaoJs3mlqDw0Vol/2HH4eeGwb
2445cLpoh7VpOOWcIVvQiiRPOz8x3loVjDv17Hh3qpZCYuGdqrEpkiTfchJNcZ2iuN8opi8oIvpk
7Gb+RHdH2I0hMpLyeYVNb1FsmB6wO7SlPwFZW0ra3xBk7E510TL6kwOTOZBp8+QsQQgEKsM+D4ex
ysMzMpWoxLXBxqCWYmYqZbcXWzYBSopBe5k/wloOgrogpr5Xpri5o/2uK1bzfFek7HVrl6MVCwYz
urQew245mKQf3yA6G/PAqViJVBq+UrYt0EAXJfXZlhCexUQJcYS4WPOwWyOZEJ7K9OT23Xw+IOrs
tESRRetsBLENB/VMUJn43VSyo3ohOn0OqCSzdJ0wzVvS3RpnjSKr1C7V0Lo6MCH5kk1+Bm/pfxPn
/l6XwMfVFiC/u+lKZSJ/C4sThQ5fD5SeRU9zM9NOmLfzSM5Le83JvUwNxkTctnskH9T5osCeUUJb
K5dIthDnnut7irrrVH9ScRQ3Afsw8DfzpNqHs9FLu9rzKB87aRG7zVPmB7I5G4bYZymiM6HGHsDo
d3fLBldXLcUvqcpWO4+FRuifW3g0ME2FaqX5U+RdozlKG3MOpnOgWKOKXc8w0j4mnK/T7CyHXbso
zr1MnzKzjCxVOYvuBLCRRHGUOC/rqAGRWLSNN6iqIvUvilnP6lPA1K2KYEWVZwDaaDaze372N2rY
r7yYn62GRtzj5fb2/Eakn/1awwOoYXiEZXQOpfx2KrY3rHYUr313FrECn3nbAoSKDbzR689/jsnl
s29CHsOl4mWFWnfOLnuexUiIzBKcy1HHVoqqUa4jGDJRY+w/BMjnFVK9zGmhzJGjijDJDLmXhA9t
XvV21hZfRcb7viqCiETi+gXTGBN1F+vb6bEVS36LP/9E8CsZN1/q77K8P+FryG41uDAdkpLOw2WE
wVeB2Fy3bL5KuRw3zW1s/64jt5/M9/GWvhkUI2aiqHfd/Iy2+YfOC5Qw4popXnqShcZqWp2sJ7+5
xX1G/cWpa7yxPEPHH9gi89nHrxoAwW7ru5022BhSNr0htB6cHGmXX3U8sci/Lgm6A4DJBQZpaSvd
q4RuX+FVgImDNg80xSXeL8KBdePnqLDd6sU2WurtKtHsIRD8j6gdpjelPi5uDulOVhxtK+verjpP
oDCLoW1UY53JEWowpsT4OLXHjkagobaupVkq7BAXWUnfCUAXs60g9fYkquCxcy3nNiJIKuEu1Rrs
V9u/SVl5wOohE6/GBHG/pAgnfmour8ltigkpcOpluRSNwnttJSzUsCkJNRTKeqdgNJQFXNLB0rTZ
Q0lg80I3ulBNRMBOILmrD5uUfKQSYw/1w+PSfZUDUb7QxU2Od9st3g2vLuRHMicu0qnyZBMkp1kH
jFFycJYPBUihSNWtw7V85tUJbMc9H4auizzffD7KDX9337b+fSon8K9OYFu9S3rKO8SBQCWz32QK
t6QSQ++1G3PeLAKbR5vXK3c+yCncNOG907Uwkg8pA/Obex9oMvqoc4WfN2aD57aUB2BJP8BDVMGe
HjgPTlEWOrOCrg0EWx1sjcxL48/9rX2cKuBmt1R01FFUimVHhF2Pc7OFK8gmrQbwTI/j+P7GdJ7h
PdX4fOy7sHWbVP0haOq3LU/kihL5aberyses9c0kVLFuvM4shpElSsHT464JxzbfCyWZDkXG2KTW
bxRdLpatId7D9lm4z3BmkFY1T46wvAJ5ma4rkkEHNYU1kDI6Tfr2nXLc+yANcX41xtfVQhyTR2+8
soL4rhJBOP8DWxOVziFk7FOajk9V4X5Lzs09rT+lWNaJWM0a4ruRs6SJpMAsgqVrCMi2LHBmrrq1
RbQUoddPzuKSM59X93yAtC6UhiVz8voACHD2GZ/Ylq4wo02w8aUE4Lb6JJ/Lq/gTSW+V8GtnbDUq
Z9CkJbSgwtw1OhIMHSjYd08FVBwkTIVY1h9DeknX+sHhRhK1BG3qyt9cywsEHkJlsfz94/FcXVK+
ikD0+ibrJlxqwXqz2DJgALOaSd+0Egt3N+V7m8uBUuJ//4CBVJrAfQMYNv4ut78ko51ppPF8Wpn/
0VyDGR0/i+dpQ4RlYXnnb6ebQObzxViNmRnrQuaKn5C/RJ8wrSSETE1SNVIUNuqnGKc76vMM+K4H
WoQSrxiRPWQn6HefdDM7Gxq3SWS8vJ7R8qDaxiNljd3yeeil36H0y7BZSbTu/njVglYPDB3zvRX4
C6fMe/HxI4UAOoG8QsBK7ZMj2Nzv0w9AbbHISDB6yJzCPZbdoNTCAX6/SpxnZCdOL6uRsgWuFafN
y+arMS+xlW6L7IwUYRBH6MeLn9cgt0oMi2XaI57kgw5di4eIOqPOH+M4N83/QHzmcNxtpNNxv0r0
fh/sAFWynvZBNp0vFl4WhQsVV/9fHnXS1Dy0sZ8ptAhrP31iG75Sg51xHmOoNpAnU3RiTSvmBp6F
1N99P/CGAnxNfzJ+JR5TqMa44YYan9lweTA6mL6mTWjzKCRwn/YxtLOfSV7tBEB8H6dif0rsVJNH
BpxxLvTDdL2y7M0WdMxY8lMqwxFj8bH/lRvnFrzcopshIZg04/Mb+iVZ+AjUX3AlebmMak0KZqqU
XV8lKmt5hByA4GysLC8kot/fc4oHI50FUJAp295/HGnu5QHIolFSnVx7Gk5iAYXwtXqfQDTnsub4
qWaFVqhmS/G7WKyHdU3riw5XE/ADijhL+bq1KXvw1q7GJtjAueL/bkEv84NBF06AapwKsI0yPESY
A9CFdlNuwPZIhR82HAZcz4P92nfJoI+TxkHisMEL3Qmn13an09WhvJQu5ivv9JUsYUICbx+GHVpb
Fqef+9Q1dMcrtHbE5iGqc7ChM8y04hPKas/RegHTdiGwu2OxpXN2aTXz1/aj/3zrOyiYYRqJP7UZ
sMkXRzhbYmZpw4GLgG63iYgyBoHIjaXPFWJAPmO4/UD2B1x9EE19o5uKUQxB+V9rgzWUNZla8FNd
O5XPIC9GqpjjxV+x/RTlSivZ9L4aC2fm9eZMYL8IvHsMrFwowdCxTt+wV9Np4wfALslzZZAitsFW
V6ltCUdymi4yDzjWN/Kzd7B47t72H2ZrG8mhcRxI0gGO3scG81mvIQI3VDIoXaMJ3OBHUUvWxqX5
QEO6a3zxEedTUEEdTSGdnGlNRVCB7jMUB7GlGFWk0Ae3JY1P+mn85NAoJS0qeNJxvv40sPxzhG0Z
FLIoyUDFIMOZVMEbPdvrQN99rqn3Ri0PZ0FKWLQ0riROOhe88YMS7L+Er2/4zrbrj01lvWPG/qT4
zPuRJFxqAYLHR026eWYPxUNIRY5ZFIs2wXPQfDx89epwCPWeTgTsYn9WWptEmh+7J1klPFDVhCS0
OXg+RUM9u9J9nfQKWpBXzEG9Yj8/PO1ti1FD+Hwe75rHKKDuQ5StqNTxPpiijxGWHj5ZWrQOuLUm
1g4dc3Y+JLH51+IlKxQSh0BJ3ixOjYAKQ/kfhM3tzZRtbiddBY9MFB4iSorvlvNzrCNJHaIO/tu6
DePrfpjuEFK4e3pPs1uOk4vZUQc7o7umXeE5Ii82N/q1N82vYmEvM4JPzzVuYfAwYELMcHDazGJT
dkXToBD97lCqM0leXouZtM/g/+9M2erg7BAYv0ASMfh+wejr7WDaq4BG9USbLivdh9MPmxAoxv7F
VH2Kwq1vtaBDLRRHbI7UutYAvOuH058hmdB4lKLSZsuvCezEcjPeOm6sk6wKTxJGgX/qQ9SF/DMO
GCAeKcFwT4P+GXTy2QaAoMaDp4kr3VxhOohgGkn1FRNluEkq2NJStnR+huH+EDHKkCJF4cjCW/tr
Jb5kA+mu3KXvIJNAxcvrBoUQL8GwPavaydI1hkluZhqIsQeCfxsmxchGA82TFSCJAVIdYobmJJjw
i0XQm25VzT2v4+yzvIT2Rd7pLZNfn4GbyPhfVlA6ltkDujJQ1WegC5KlBvjBf1uSB9z4PgZYh0r/
+CGIDmP4mcRt0CPK8jRN/C8gg+Jxu6jJEKQzvUXZXws2OgZqxwMGX30bwYP4goMtx8kytIn5IMNs
3Uy3V41ME9oc1tJi7iJPB9Guspo/6F1NmrOvOC7JC+Pia6+Fu/lzbQSQ7xMSuHCNqbw7U2o2liZb
VRX0LBGzUR4UytRItPMwfN7qHV7uO8BetQQ6woJacEzwPvFS0NdPlQ51YJIvYab/isJS5Q46/uKJ
IRUciQ3RRa7QeqmuVHlZvf0LYGUPFMejFPNIl8YcYxum6Lq0G8scE2aLy52WKgJ6GreCnfjziL9Y
MSO1rxRUGm+ziW8pRdYFA7waY42hNrkgbtZi96HAjstgo5goUyLnnY6H0gF38krLipEcSpMA44UN
9gOyg+nd5uBPHPVUa7GdV0efQVobucfVDchqH3AM7nhtIkA3FWh5DKgMBj+bsZrgrRqiNP1omodY
B5Ww1d+4KZbZKvdIA/8NV2eMRO9UU9krdrapSE5hGu4GDNhqsCCDd4u5uTXZpu/K0cf00ZGYOOdx
h1s3u4XakNGCRJCXJHemyr+nHE0pFCeNXVlwi+F6sxvKZWmkwHq6qjinlFEdZMCaoE/8oYrCIT9N
A2Qi18T1KQ/uS+bEuxy+3uf6S/7mQ6dl3FUEwAbyBzQeSzhT/OvyX5Td/3bnbKmKFeooLjWgHjcI
kx7hse5lA4boAfIOBZtDnqeFa1Z4b+E4Nvaf/W7d003AbvO0D1PTT3PVTD76U4b9CYv0QFhPrOyt
LVOR1/cjKGxiXcf95PxA4muINFzy0qDDno9cWnb/hadJj1iduZyOPyOYUdgw6a7Ar+kC75hCK222
APkvJDVnPkgus94JvUe2V/82ZrUvKdF2fdVkQ4y0MUbAZibfdJAFD09TQuCSUXXCD9La3wjZKfQx
4wTyFU6E/qxKI/U6TzaIJRn6ULx6C4Dg9Rjd8+to+61g6BIv3mi+BJzbFaqdG09LJpgu+hkB3B8P
BCqY/Ru3+wRMLh5zcxfMGjG2iHJsqzpQGPzlMQg+ilPirNh+3Ed298aiK49xVU0dHgAArntzqBeL
BaVyOtKrLS/yXVNYBgV4TcWBQjDfZpMne1yeZEKFscstiatzDutol52DR0SV4691g+iMa5Q/v7WJ
VQ5bJb4YlFd9ENNnyym5Z/bhsWdwfGLBjQXxDjtESLax1Wmnje3f93Jqw6EuBn/H6guslBGxYaQE
WLia0yMRL2EyPZS6B6fBNBjxprMA2rC52fV0GskZix5XyOz4Q12HaIEgvQHEVO8hbfmjC/prS8hQ
Tjh3205VqeV2eSixaGS6WvSFlQ4yBiKGJO602OIGAY0MnlhJuaqnwlEawW9S/8UHJEIFWh422nUQ
yfk/ol7EyV+MhJKWaXu2hHlXk8kwZg2RNLe/oKkcCeaL92TQR+DUG48mDyVSSlm8TAkws/NbeQD3
oZ8O3wg5gituBsi4aANXG/rYwvFQHB0PUR0WQ8oMBqp4lH1hVLcbrto3UHA7KuaRlz3YYkA9iqPm
TVKPKuDFI3QroRGsEWd1UVeX39gUvK3bjnyFrc7VhA1nVvmMMa9MHNLDAIlR2F8w1VGzN6+uX/tA
j7DonnY2pEhPrbli4hkbiZ18Bql33dNuxUwUXzOK+0yda64vvw0FkgnuPpuMMD6KPmP9W3W71xh+
Qkqte0vzNxoqDMp0f/JKRK+oM0ysmLD6S47tVBXF1oUkXJQvljNxBrYhPzl6Vd6awUPzizzerqEN
HytLy+ej9p6ZOYGnEPcMZifSoeOSGMYLx6f3I85qDQ4yAmLs+7m3TeqrtteB/UdXMX6Vl7jJ5mrh
oacmKbiZJoR7fO620GZWkTrLQVVchsRY0Vrxle58c35ZvPwWwM3nF5ydwgGQxyrva+/+W5EyVMP0
2QD5TokXk0yxGa3GCIfpVHI87cEQNBEx6ukh2Y15QTQYlAQ4AKxA4wsvjDbvuR9XP+31tLQq3En2
mk/TpBpm2COE07V2Tm0PGkwunCQhh+MTARKkOQ4lr2hnHPZWVrMfchjc5rA9IFkaMSp0lgbEap4V
H4Eh6+m2doDWRSndzuojZGl08eH7kqUwbgAYpZIamh3++fgSZkOYXWhIFfw2SK2P1HHZnhIAfngT
lRVfRBZPRmz5jNxM+bgIpTdWsB1XZw2z3c21GExtzTRZmQci7nmMb/D4jthUsN7iov6eKLCvYP2g
Ri09Hi7kw/OQ38W6+2Om9uGgzAxMWiRwF+zv2M6boU9B1yIEG5tWswxDOc2diegsvN+YAV90wbfh
iumGiQ86G8qAgCdPpBaIqu+hxMDypqCoCJtC4jC3kXNcwx5EaGIZz4DnrI1/N1qq58r1YLNTVAoT
n7Vm68wdN/WiHQopDeFPBkBGgn98kvXyBf0SUstfLsCcTg+tJW2LJRI+hduxvSEvp8VB87Sv0e6x
7Yi6wMPOaPCundPWPnT2cM/Cx1R+ET83ZTuplqWgKiNftovV8hlc8pzPkqVSKlMOhgNWff6d5fif
tQ4fmKa+hu/wYrDbLp4SXcttZJYw7RHCecpNvBgGY1ceaD3nFdTrvJZcuQ2Ocmw9WrGAoQ/Njd6W
g97tXMgle19ppjBgZepE62sEy9rgxd6+H+TYhfg++x941Ajy7e9xszdirn+KlwTk7Qy2f6+QOrCq
kROeC4pT0nzYQ5yJfmU31tAPxhIGC37FrZYB90FJu5T8o6Yw69PUej6mnjbeejg4AyRaXgicY32h
Ie7XrCvnT3REUTPwu8FAZ39GjMmvv0sXFWYFmAzCxBPV76W4z9xFfngpJKPk5jnob45T+BxOXLJ8
WxNDEypZtwrGpzam9dSrxyGh1G6Ji25ohNcSJif3WI6Sm/4Ux2fnSInGTWHESmll2oZgW6Ttf07Y
wIWD6RYJ0475Y0NnHahL7F2ZLw9JtUrl8kSJgMdoWP6CAPqyNA/T4go3EIRid4kEE/AKjgs8Lquc
XNMsklFj28kHW2AUAEswhZ3ousa8x45CNt4GOrkOLauKB/WwJVQ0SZoalgZ90TjfdqGJE3dhD6cY
rFLyeX9F41GKNPO7WACSbyzZCPY0BLTvB6rJKeHNE0SET9+uX33RW5Lmc/dfynO1RsATrk/ZK7TM
lhq5dPv+Vz8riHNYFzeRmvUDSiGbHQ+sObQmtXQrwWsUYN5TmMuf4QF20f/MIg7QkCT59/z18D9n
+Td8nI9YA4jB7Q0+212mICu9Jm+KRykyvkiJfpV9CJ6j/ABdtOHKTHCafAraUgVAbIxdMPL/OtMo
cwOQI1A/9mt4DofOgbJEgFzICr3HiXSELh+UCHlaThsj1xkhJXHP5+W/v5kNsmpSk1JKmxt7n6Po
1nuM3kzIu0ByhpuZZj5+Q+sEeAihmPRj6TlaFWb5M7f4D9g2sGu0Nn3KoPBdVmj1UzRdMB5rXnLR
z5tUhu2HXld/7CNwSquT47J3Wq653NmTMAYlsNujAwAQ0DNgfbgMyU4gSQsoP8oxbDGyQFAbNcmQ
eqWKWQ+kd152h84e16xOhxQ3SJnH+cL7bsyJilARvGG58ZVq5CXfEPazzgdxmnmMFZ9Na22AJ+29
a9Bvif7oG5xt1uIJcvdzxRi/GoKQ0aSIy8h3CS6xC+bRWRw81ZhXGjsYdd1iPLx2m/q+P+fLXVjw
BHK/voufshvg6sCkXEkJAyFF4VyEbaf4uWL20Guc0Ee2JIP3ev5kKzKgTm4PvOK6zz16gEll0loc
4Ju9fiWqH7hB44j/eUKD+tVEbeYTkE4S9pAqcfQ+hTSv70iTOLwfd7iWvqCVaBYVr5k/RUOxWtmQ
f+woMQWikR/leXIbkrTz7YTQ0ymUtMQFQpZ6Wu8uXDfLcNY73Vasb7aMgewEi3OnnFBu4NNSxeZq
acOJeDBPCbgwWF1bu7INNum1QPaELawl3Azb6Rpb+MB37xIA0sR4aw1ksrgsvJ6fqA/RBiZZf1d7
YZbcBoXtuLzf3vWLlG6xXpEmUPPl2rsbwApk4lyoY55geHuQgGG4I9NNihEjU/UWvEX6zNl8Q0PK
g5qWpVoBMwywJaQKXJuvBX31DsKmHjArrqE0cKeOxnAChIxMMH1sPd7we2XUy3eLmjhuv0wiaD9p
O8xWHIuYlepO04m7C1Te3aG0ecG5EHhm+G3yqZqxNOUmfkAW49ET7oLt4NZUC90ql1xyk0Re3EKV
XViD+pwSMBKuzldx/vkRZfY6y8Ek3k8u0hzvQXOOReknwk91c8+Yawx31emIKtI7tP2gwXJRp1LN
/aQh1VuIhHPN80EAZA97xoCxA1tG4185Q160sQ0Lgr8+ZJjEJk6IbY92DtvbeULHY178nfW+gq+y
aG2hoGRsHWfJmdTaJKTHafcT8ltWV8u0Qs8OSur3ph1w4UqAKWM9kYuBALfcUNyA01+Ts5vNNC3f
t8otI+/gFmjLupiJOqr4BNAJUQnm7NYa6osESqdh54CYJ09y43g33EXRBKQE138KJXVEQ1lnCTW1
+/rx0nGv/jUxieqA9HAAIPXofV0Pdzc57Tj5aQMlkeyN8vQT5EW+3+mQENyhN9Pe9VJhzS7dekFe
nkU8dOaC3ai1/XVj+9bfHwkc7iviCC2f5w0Cfe+a2BxFde+7Leg61Yhg0EUpwtKTd1QuEgIOvKFp
ORmIC4NUoA/me9SQpZARdmSKtfpYN+Tj8hpVM2qhYbFfUhqp4OGgm3JbjHV5azfhdpe/FsapiEmB
6GM62SBmoK/+dNj1vAmCxdVuG0LNumwCffsU2Rl0hb26BCy/VoAbxj4IpboRMG9ZcuOa3g/x32bK
poHiBrTcNbG/jn+6KhVKR3PQsDFwjQNszHkIHvk/+fRhFJhEKVADuIp1zBHjxf7BWNBIAEXyDgu7
Wdi6B9jIKG6UxJvEp6qmstHuBTejOox9pY1QDBGlnSPH8EtVeUezT7RaQcOJw4d+SeWS7PQ67iys
4eQTTsbLecCoZSmIiZeVhipf09nPrcJYbXG3uFPMaIApyJiGZ7XWgLtf5R5ieMFJ87WYqBn2h9hE
xvQkWB4XWsvnU+lpirX/Ow/GUbI7ZnhnB1LVI55dOqvEWTWDwtGv3GB1Jvb+Ti2hv/GSshKn/Sal
d3eRI8ZXBe80ptJwh3KdibD/cqULlZCdbXVqtvnbDAf0gPV+Oz7yBPuAhaeUBGPsYYspEADmR94R
h8m4QHUMtZp+sCAZGlEUJyiCmOiMHJrKCxvgp8LpK0nPdQpfA4ZJcUyq+aA4B/sjAzwyaGmsE4uC
lP5yagGpcYCFzMHyIoDRjdCE8a4VC81lZM7oj7nUaVgtDwCFIwtuQDujlMdiD01PjF49ugrWQU5N
gy8vEKAfoFtWF3m1DPYkmco7BcPzTnE742dpulxWaWHgBCu548oJ0cuRxUX55MW7PxUsJHzM8UNY
YkMkrNTDf9QFOIJBjwu3tfEKGwQGzBDzuwwEmYcCo7EtMSgHQ3DVeGy4myw8Tc8SPv/e7Om2xfjh
Q7vL+oNZa/LrY9yTmRrPjqatkJCDXqo/mPODRWpb90u63Topx1+eKpfVdS5wN063bQazfOIIcb7x
I3ZRYSRrCWO6L+KmaM2/pw8RDl/3Qelbz+3hLpSBPsvKq2itxsIc7pS2/mXVO3hTdYUYKZzqtZjV
21jo5vUCVkivMkyRUcjr2xAS1boVRB8/WbA5CmlBKgjz/7n3IV9ijFVpfUqFFO535JDIxVdm3dp3
j3cw9us9TG1jkIKxtxmKYRLLpxpNzr2yuQoFXFTlUCs6miJEgCjb3JWMbZr1kZSONLkeoWHFC4hd
n0oV3jqbw4HN3TQz/6VkN6a7byPjvlAkOBhlSnc1Be+oc75DFqIYdoksUDJNakO/mL660CPeUpLl
xzX2SZhb34kuQyMMm7jTN7LjcpXzxk6+80AbSRTBqt+rT/aRQqtqEZeWgSOK8qoFv9mlzNd+lWHQ
+u7siD/mAeTCSJlfs+MZ4mMw6I3W1DyzP8EbR15nuqnu3nbT+Yf/P9pyc3oRHkAy2jWeN/Jcw1fT
eBRsDwKG3/xqJ0OdjFz6NeVGAqKXbxjXNWlNfTYK5nUiRJe5wpamIydLAOll/oCgd+wGn0N9TW+R
WcMfeYKdwvFuw9MuLbVrwZA1cnmYhWSVZ7g7ftYJn9If8cCQuaM9IzwAJBtXWjsqBPaY6knQGZri
eM1dElk/M13HKVslnlkNbAqLvf5zfaf3brpoeP5vkCNERgiFMRVSZskQMoltxYzku+4XTtEgtT1R
3nDl9iFL5Tf1RhtKK28mUZr3nOKXCzkCEKAiW3J63Pdi6vaQ+SyWV77PAcdP+OtnjgBSonpj2A1Y
JYGpBW4O2LnYxKEqIiD8GyHukgKZLkHRY76VlvFqc75FvQSagakA5dF9R0fanaGMEM3qVpp/MF/r
HKBF8woeNcizHuumFQetZu650jcbbjEVUxBJeOjK89Z9ByXMCNRxQsIPtuDxoL6bireT7wv1yt/O
WBeeHhNb+PIwW3uHU4jeNiq2XQA4q7YgnVt+GtytIRod2pA+7Ep8F1yNj/CtpK5Cqa+dBNOnwMQO
ETReMPCsOTio/69X0r+DgH5QsTRK1BT9VMpuxmHTPQTRr1SGpniKn2uvmONRN8L1uSWAjb3z1pFS
vpt3VQietgpxGZmZwc+Fhv/ZYPPujqIJDKImiT274xkyctzA7I1ApUeqw7MTv0wRfZrEL5cmY6t+
Jt8hd6ZCIrIRNJjZ3nx3bJSiCZPhAwabneVxPCWZHc4NywiflgYp5RjWoJ7S96Mp0tos2guernry
xmKGkNJcIuToZNgM3778AqwCONnW4ZY4d+UEB/pFB+O8CWUicLs7G9U1dRF8Mf81en+OgFS/qfJB
6j+5s8JAcmxSuwev5OXhAP5m4uiMOLuSisTxgF+sUpo4iwGJIYd3x6zBeDj1TsI5dM4zHYrBhb6b
2qvZk2CJ+1FUm/OgL7Rl/WQ18/AnIzkGFCzqkN9MUtexzXFv3+c8Eqqj4IjAXwPvUTKXwAknEoOo
S2ki+4Bq4MF+elE/T3qioeML2KRJFD6dbeSSfp2iuRgGRyQWJo+CkRP2WWYHw2poF1OdZg79HI1h
5fngG1KghUoTSR32tk7MYTj1pDRV6nSLddnX/VudpKt9q+3SQzLqr3pYeg14JTBoXiH3JnqOcf6E
xX9qRXE2/UZbdKorxR3qk3IYYtph4N/p2TNWqkGAqglItR5/coQWxuzkEa1YOLWT5pkAibfx3tfb
RmIGVBiEFZR6ca+gOHiUxExfU+93ES6yabW4CO/PpgJkbZdI23j8LPAhce8+IBU/aGhVNbcUH4EA
oyl49WWxIyMFowwg6tqnmhIVHGaIHmWKtVRBakavBSKOX1Tnr/BOUM69PQ7zIPwNQkzW2bCY30sf
+FOzaaOUl8SV5lV7bTbEHPYJjlgd82sIYd2mSfN2nnzByDUnpft2Xc/S9Q5pdW9AB76bEhr0L8sM
VXDXvbQgjNFXKrdYGOX5pNKOlN5oxhfVGlzW79HDwyiyA5GD2G2UGU6TXpCYCksONjTshC7ksmxo
HE2lxffsZF1yK+G7be1g9yHqyMe3qHtDs8q4Vml0tsHdHgXCO1aGZG8aHDe7z4oL4kwrJQICNyIt
3b9uuA/ybvy8T5wJg4Z/qz03umT8GT2mVm+Rig8jsohlvItX8/ItjkOS/8MuaQSUbbnzQG7SDgH0
wfR8RVTwG6rcIQMRSzD8hQ+4Ytv9lpURP/d+DNA9MuFaBedaUx6Kevyz1tD+ZP0x+42SohUX+9oH
kfEkJa1mGQ5daIA4czyIcAAOWeWNrz2yPiD+eNUhy8nDywBGnjrmojJWAWCB6HP8RYMzysyX3wod
8UTxjlJmOHGHxzr9zWb6YBf7zSUdMyED94AWshvHxd8czojOaWrKYfW0/WvQ0uovMXtUGuiu63Zj
90jpLkhhwQkijC1reob/SlsNywM2uo5MyacoPHZNUkldKyGQIiWvvSYw7IbxXGVJdEHMQnDYikus
YSBn3Kv1Jbz77pcy8h9Yc7CvJDZ2vqbWMm5DcpcBuJQPvkFXicdn35WNMxey/MOfj49MviNOKAd1
aP+gqCY+SztlI/1krO1tge5JHbT8766COYPpuTWj8x12F6Mr/8vRzTtvya+VzCTH/tooO3Oy2SmF
wxXL3vgC8M4U2dvFfNmK9YuuKF5QtIQfbOeSOSM8VVq6YFuNsCd1R+01xYR9skkbtq/dSBCpSu0/
4FAZ4jQlRB0fhsGP5b8kKezWIWowYHRxry/HHjVD/oJSOIfI8VrdLx0F1DNALrc2+2zd99TQ6UoS
XLtxfebvWHqITRUIsHh0JcM3OML06sxu/Jnc1X/B5fUWO6d6ByEa5GXVJfvO7w30b/AXFEZlycyf
nxJVr2aWlZMk+2XcEqA9c8pnKV6u08DGwXfYcvVDF1A9PACmpnQb0uH1e8SMoKI90b+w3QCU4PZ3
7Ll6QYGEZzk4KypLcbMt6tkVqvE2mZT0xciachZuGT8greuuI3sNu83WHaQZ6OGKjxf935t2aIeK
FFN5Z8RWt27sPaUgdvaDpDgNPHFM3+/kQlSZPg6IRhqiWVggEA0lxoFZbE3azS6PHIEDERX0C5Z1
jHLdbWPcM62sH9wVoKFXPr3AbmXa1dbjX1aI9EoRk8bE7FlFQX4hAIpjg/b0uAmeTcJC5R0OeocQ
CvRnURoMPMJE/eJQJ0u0GVeJ02Zca2pOvoVU2KoZ1jkmBqPz5DEcIa7G2qGqhb9oF7fv7Np8xdkt
mAErYpW9QfiCN33R9xRWV2EJ4CE8hox2RQVHszbbwW6MBGDR9oaCNyzcmuY2Ri787ToQw2A84tIY
o1TmQJ7rjkYZEbXMCVa35jBoHRDaLdYFVK7PJBHNwakR6/9Ip0Kd8FTG3DOJNhfBP9CYs7A9x/kb
lx1lMXCYo7HWPODU5Wv2nBMiCJFnpAiRvy5RYwourOj67veipPFQSPnhmAyvGgEB8lw3ydfQbDXF
DCQ06kDaX8RpPUwzNxJkkhPio64qEsaq51XEQHq4qh3WoAnjAzWclyRiFZVFHMdzfCFqG+cakYea
iXjZejHAzV/cd6szM9zsgqceQGeU/9Hb1sMduhO6luV6JTvH6r6AqgxLjJSHK3iGU0Vbvv44JFy4
uMX3F3BPgbp1ZTrTINb99JbiNNe0Ynhvtc795sXDLVkUyPk9ApucpXIJocEONGd7dXlr/xThfNAz
7vysV3FyT6F2A5+LGeRfeKh2UCwF2ZJsMjLMW9F92wgth8mMvV+H4ipdD8ixs1doXw89gKuFrSII
Yawphg5LEknhV42voi9sfYkI6VI/HIIXFI8FWlz6XvmM2LLQpdZNwuo4lxp/Rwoghs+6DLphQsBE
/b7u9iBQm7TLc774w1hPXISQQtrAANZ2PDfAkm8i0jEYbxoRBTuhT7HZl4qDDCyJiDI0lizBK9T6
l3AWse8+YMAKhOcBCaNCaZW5UCJV0WJ7MLDZSv+3GVEJKgaRrk75BQbF5U+ohH4EENAXios0V+5D
Rmqlhy4KddqaXNtCkWT9JxOQwaeUKC6U1SfHWdTnOBLgMMcnjrDhlk4Nd2/fEl7xTCz+WDyTx3+G
aC0DqBlOerMF9ZqHUvaVJkYXJxL40xGh2HuFQYW9W5m5tcoKZA58aMqEGW7lfccQmGyRlefh8H3V
DzsZyKhaS/NdzEEoD8KB5ZYpmsxcYphQwnVk/RUq/QFXvL9FlEfotipp4c+M1n0X+ypJW04RRRrM
sLWQRENnN0LLoaoW9DUfS/dYXtsDWVCQdUAq5RrzOLGMSxyw5lJ4L7gv94qytYn/bSKFDJauFYPK
Rc2Y9rLQbD49MCHJgX0NBYevLsYgqdphwbWGjY4WczlL27a+mL3kmcH/2o4upLd5oeBcpRRScmJ6
8yfH1vKq5N3DArLjFQT2Cr+zjL8fcwMGRGvdIUjQpOoMB2Z3SADvJcYYp8Sgze/YwOpFS/67Oe7q
lQuJybbdUOreGFRbwrjgxpsW52NU+Dan8xGPSXN39ZjufSCJlKSKwuQprqIFW9lCjrtUm8xLc68v
MSB82mAcUqJ1Q/GNS256fv8DJaLR2/ljrRkAspTd245txSbej4HbCMtWXAjkkABYP0TrfxaIrFrD
xZ8aJ2+UF6+nbZh64Gl4OOngVThzqQ7zqSTRGl0d7xGblU5jfDqASrYez2lKl9+B+ujRi7bTi2Kg
OMJIZV8MxpDUvmM/T6n0lIg53KOLZ0KkHWcgS3/ndYiqJbNgbtX+Kr0XineiatPDRalQQlurBNZR
o/CQzskj5HAI6Px4IwnVgXjDdTzC/XwUgoduOy5BbkOyg3LLBHJ/pKLOKNsMNwJJqrnXoVCbZAhd
IHj6HL8WTk+475bij57hTlel2zeDCS1FuHxlTth5UBOwasYFtOBSmjtx1mN/9w1WOJadXe6w8/HZ
9SiGJ9eTYT96Z/VLShdvaMTZQwPmtJZWTJkt0f1fqyPUEI2N7MiEeAB/JnTrONV3Uc+qyRR9gVR3
vVXphNuXaWeXboQBdkKiqc8fk2lodHuEHodmJ/romfDG3YCZZ7nfRAjN4F+RPQelr1HYy5pHaSrl
IRgBeGYBHxE1OUOCwFL2UCx0KMUIZj5ChyV9bX7j+UVSJ5AB5Nu+vqYs0j7+GV3D4y53ZcRKP9Ra
2mvKTxDek7OUqE+28nItkQqXAy0hmLEtoDpp5D4YgFeNfULTr8T2fvQ62AceJgr9++fB8nIaYfSQ
XhoFLsRgQt/90UwxPiKRV6/8TJQ1K9+E5f/5wuU74EPYYX2qDwtCgTk4JnsfUl7kEmiJ1yBnACXX
rcrgPGSCrqQaMr56ZSR4UbhkCxL8Ipxfq/dNmfHx2cjn+7mIV1F+DJXC8bfVPILW4SbSUwEb7fCl
t69BV9KR6zKadv1iIgxQZLfWCABIKLUxErbhsliG4zj8nGBJrLupY8wP+W2OCwyTvtHbJZIsPbOa
3yZmX1g74R9OozM6hU1+tNCmwe1IQLTZt7j1HUwT3kIyrapDFMs/4CORHZov5WiX4mRrvSRUobWV
5C1rqTIbaL71Z0zEVLCtoOPr79udHRe/9WSAR2y1q2yjAflUONiKyy4wskmaxfi4QLWmwPlyZ3ve
F5GZKAaiJqPPGo6FY+cM/c9CdKGrnZLIThK7PVU+3CDFSJiTMqPfTYe0SvHYJB17c2q2nSAnvKjW
8C98EoxuPUMzdUsPqqwXc0QS66Yl/0c+13Zkf2yJt8iovho4WbzfGOzNBu3jiwpmC0F4eUyEzgvA
xPpnkbXl98zd5EbV2I/qtp6a2yKjimelwWplCoqKNNrYdfNNNfvbqpT5OV5/MQpE6vNUjzNCCHia
Qc25bYmOwA/E9HgcVbouqN+kdui0phVULcHA+MrL5SHQNWvCunXykGYQwZfkKAF299KZMot8TWzz
SBEU4v1KU26+3+6dNtSEnbyCtyul3Qp+FLg3DvxuD8Kc7g0xcIFSibtLDWq/5n5OGlxh6dh4cyUF
rN3ICh7KLGcNax2/zGSuqP6RXgKSMc28MZPT1GRCQsFFle5fSb0nGjdnYczzpguwOpH3lmqvWl/P
ZCSnSDvFBwAkFE5W8pYBbJlbh8belXEdAMVAfKEbFmhPW2Dg5/1eiy8kM1Oy/jGB5Xc6zT91PGXi
DVrh+4bIO0XX/fbR3ch2l7qAGOEpdgJJx4Y6dw8e1vnWhqUqIN4yltRC1TnmkjQpPCpDohYbA7MN
Et4HsiTUUziQCnfdIWIGZJDWY2HQzmIjrvmNnKWXadH/R7YN6ehvxXJ3z35tNSJWBjMO4UEx5Rup
wxpR7qunx3HMFS/RWMCOoxcLvBcyzEcoZGl3XVXE2rXiVW8i/Sw01K4Usu+kPjetQpb7ddAFN+oR
OH1wpVyZAq0sesfyVFKm5Vzp4QMwUzQ/PKckNWoKvaEjOeue92jFKEiH6qBioUy0npNArYh/esOF
+qXBnq5Uc/MuGkhaEynVweEPUPf/maLdalREA5IVD1q5TdV77STBAJ/zxsIRyRqEQ0n75H3GkUZI
lH392aTkRyba/A2U6YfOEuBUKl9WdSrVk1KS7zcJMC1BmLPkw6a1CMkEGUffiNxrpQ+iEtgxOiN8
Pvcxp+K3GkfTr07UvhWhdO9OMmlcBc9Er4FH96GRfYoDl7bXOi4vOEv0yoaVcSssABLNo9R6c1Op
wvMxFZRfka+1dVYl8bptesned//jLa1nbIpn8NXfxh+cTpJssWn4iEqZSo3CrheZHFMnaqzwawTg
6kjkhaSJt3mFHYMNoNOaq8ELQyKknJBeBiTa1n/BqDnCJffLmu+z8znu+csRd0YGkvJDnA/a4bnj
dwbyDAGBs0N3M9YlMUCtjtJNcC+00/3DS5jcBkODGrhsx68Zdg0ZlBlZWh4uAklMI1vIhZoj/5jF
vRIj6PFTqnSH3SSacooc5lFXSCD/9Q0Cgo7Ot6ioq7iiJx30G4MLfrdvomVW0zXPHbIN4bthsdLo
TlfrPeQK2J/PppCeOR8KKLMITi6JCtS454l3z7KW6Ok/FNL7WF3ARBK293oewHQ5nZigZ6PKO2VQ
5x/2hi8KYIqoZHDiD1LVzIrfy6NFSx8o5fpEmJJdkP3jIzEmMMR3w7SVwEZ4TEtKWc+kUZOp6h9f
yI3t52fkV3be166Ef3FVMbIjkP26JfA190oCQx/JAcf/lSUmj9Bz6a6rpJm2GXwbn9iPgQdAI1F1
3E4VLpc9ZDUyWHxoRfjYqZuChQ++0gl8CCU7L6msdxIkyF5aK7rEW1H8Hk3eONYeS4M6jN0FFTj3
Mp80Za36rznlhTOQ3VI4qDYwPdHKQ9A7NYer9Cth1YyEQ1fynfY4bSxHiJmQxhuFbGE4SZAoh9f1
qrs9kfysMnuZVE3WVVwtI0XzJu+v13ROPxT/op8uq+hNBzFWxkBwkb6gQ+ySKCA11OBZSc/T+l2h
we1KY0eSZ5Um25Tybt+QgFLIa5RpdxZ4IygA0CCI25zVrq+DcbpiOhOcuVMNJZUKaKmzozfUhRTT
+GS8Aok3/yYu6HeKNCnKtEUm4DA2MngTdmu2sM+CsDCeyk6VX0cdeEi0LUKL69sIBPWJw6eEGVf3
grD+QUpwEFOkGxl7Own66VE5S5dMY5VwDnBWKROFvxV5XsWJFhcvCxDLJGBgS91fNnKMH689fPXh
k4MrO3oNt82Y9D2uhcXhkf8CjosFuuhCXZJGUve/hWkv5+FruviZSv3SE2f3+pX1azYasmaBXxEr
7CPmu4Qlt4aAgf9RSpJDH0nXZlaB1v5t22LQkUMNJS55fU7VHjt/68Fw1PXyPuMyHg2212hZs/Gk
Zbs+YAxuXBZX6cd/c7GfhgUXOwkY3Sd/nmDogtbo1iEQM1TpOYtojsWvH+sYDcgVJKgj6zN3ALv1
wH6I5E/MZV3fRm9nGs1ajB7PAvGnBeHoWnrTL1a56HYyTPxpT53OjKX7m+nQz71bN1LLYtWi22E3
rEAWwSuGUUDhV+EaVtbCvciXOGdUK9CRdkgTglwtSVi+FFb5LniN9Vghs2MaBDSMfXwohznyJckM
5Ox3nu8ugcPX0yIjYrXHl7ZcxC66h8f1/SJPU/TIlC5Awt00FjUz1LLkBuQNPfLQkmATujP/XVMc
rz+dEJuTRmhs4mm6yd6hwMQhwPKBGq/6cb1bD/7rriMn/2p/CTlPeoIp72VHWiORNv3Mbyy7rbBY
b4GDa1Gh68+atLd/emcHV4z1Fv2KOZEFy/GX3bGMw00Id2vNEgM0YthoLE3mswDBqMS4JIDTdxh6
LvjoavTHc9K8luIxZqeuB5X7GJOPJO4HOk4rS60owvvcAWZrWa6MrIiiNGt2wBlqgyLNJHnv/VgS
WRA4iUHZn6n1IdCKQ/wwj7mJTVoWosEqUNbi545pWxpX9w2abSrMiFhGuuzTzWh7jGjYskiienCj
dmdl76SNIYEwjpoqffnPzUWjVaJR/6alJ8cUCngAYaJAnhdI1yo3EbeZBp/iv3xSbczpU0+vmNce
sBXOP7J3OPtnabdKBL/GTixAiA7DcpkkHWgyDhfxO4vtjvSHlqLNW9mIv8bueoF7hrNbZl4lXt22
P2banWaw4wQ3QK4Cb7ynNeycfrWYSI8gmXMPl7gzZ23DgrjIVfHp1PoVjPb2WPWukZ/MLzJXML8m
GSjJ2bEp5msTmDM8Zc2giYvAz0/8w4O4og5pnocRifgli213+/tkS5ROMLVi8uoaSotDKNjDyxqZ
JjReN9HjinjQ1aucsW/mloaROGCFtxqQgiUAC5VljMH1O213sT/3dbTmeFhZOjdx4RxvLBdVESXC
rv4pPgPXwaCHI4jWeIFN2dwzB5IWj0HLsuEaxGe9p6JvrnAbnzzn8U9QxBBiWuv5dwOZRwhgV90K
zWdKnWnkFaU0VWZx4xZpPfbLKxS+Fv3urC0loZ5A8vn5rq1w1fFUc0vGLPsfiMQxb2GqrLN4Atmq
nwOVGHtta/YsVTd1hUM0Csedfy3ANyioxOMYgAN/MsqtwS5O3givCshoQ7ZdruyxIrFHHItjmIWi
eZJrhOEmzTeQqYByh8osFLLma7lTbJgUAVqXqJb5GEbgCr1/HSzoOAwH1qbW5ymXxC1r2ZMuFKvZ
wDqttWGNwxUaNunIGdACoWLJY3xJFFGCdITxRwRn2dz7Rczdf0qei6RMMblFUO2V4giLvvSh1DS/
t49uo1RoZ1qS8km3ZYvp3QRBpw4jd1j50IbtjcwNHCy4mdOGbtfgY5PWU/BuQ5LJBHWXN/L9jnGh
dBQViwOhZFg44cvWqGlvE49pzy7DbQ+T7r90CmRdNrmUuXsUwDT9JJBVFjah0TeGWafPi2Toq40g
Yi5zG20EYXsXkAUoZj2SBeTE6d1heUSTYotL50c5dwVRnDFRHI23iY1OjCzFIpVa7KCdGVSQq2Je
GY5A5Locg/izL5Q96qu3t0VtBK8eoDZ+KzAiQzdjLzpqMA+b7AKodwwV3HWw3UZhdTfCPNqIogxv
ur9rQJBTQF/iYlwOWOpj6OT85rP1a/oFlM7dcBjGQmweuMEndkXEFgHmgENwb0abX8f2AOuqH/yM
vJMNnUo7gbhUjGgzFnAJ6NGSOq28d4W9+yQuUtmRXhZiqCePUHIPPSkc2pY4vgW0T1uE0nzLNDix
eVukk0doHXGN8vcLq1kfP6kRabp4saSueYoHhRhsBPCWqWm23xENsIH1BpZq1AWS973nVEk1vfxW
OHdsiqVl1SpbO++216oGPmAEMW6u2EMbELpgu2+8W/otQMUU8IHyPrHeRb8hjFIU0Mge0Buvuqc0
bWpj+0cB6AGGwsJ4Ji8nR9Rb4E2lTriUDKDt0S1WEQa3gtfexNoK62F456e89kcQi9ye2woQQk8D
+NIPgDC/i5eW30Rl7slDio4pswoIvmEtQeoa6cP/lJQYLwoqnNWNbJrkfgGq8ucdmBedf51aYC7R
pdtGbGttw2EsiN07/Lz+SafE5ZgU6SbaEVH9bm3F1u+XeMQfinDhVQvCblYEJ+0Ks4ZkiFKFXm5p
oQomWVA8dMZ2byHW4x8Nua1cpA1L0ZkSTLztxJN4uaY7xrIujPg1jEkQTDyf08tK9v60R9dZsI6z
IX9UzF+FZhKdKUN4B8U4E06pQ0uUPsKqwck8RvBI0+dkNPs1nyq00CxT8n9WhbSqgi03j7GMlh2+
BuuK5SuIOty5o2wZcEZ0r5xqbWGOYERaHAKoZs2+Y6Z5rRrxtX7sIdxi1kvtnxFIV8eH74DsfKHn
CGDI3y9g3T9zRaRcKWR4mUyYx0EawGls7+kTX2oNiLCZn2FhavaAdp/85GLiN9Cev+oJjOSpyAvZ
j0MBB3lq+ZGQOFAN+DXGFcn28tiDiQqFtG/nbYEp3WMKr0sn1NGs7sSX+b5AAc2odM5kmsTHOBgK
9cegaKySK1hNQtkkmL6mMM/UtWIUTJ5NupQZVHaVGuezwBz1ZdA0hRVjolLWpWjb9kmCS34RPRhh
KNGugor+zaQsRDBFu7wbE7wsnPCE2f92cFgOSJgatoFptwSklMjnCfikhRLJs+MCsJXm6YqB5+yY
BeRz3GjFObm6yxSQCf9u37jPzu5HHWFUQyQOGbNzLdzXvVlEe/4jbCo9j1KbbG5MPDWG9cTBtCnG
LXaYudNamvP0B/fFwFTwlD2csdoz1X3BR1HXWJ0/LFfit5hQ2L0zLPT1VlI1Z6um7GVZyfKgI6Nt
n6t/pNRwYUncfkLJqn9Sd8hoI2BTsIpn/VT0XRFsrRlwrPKOnPpgLuYdf6z+BXj4ZXwEyESKveDO
HZjPXDexsNAsdJwfBYAL3u4oY7cz7P6VSNNhL3NdKp1pZvk8aViYPqm2yK8e9Gq83XLhDeAfCYuC
k8+JR8ucKBQchx9GHSRXHBwWBu1Sx1GGycAiDqLg1dvdHT7VeZMW2akhNH9KOhQi/eh6luS4ZFFJ
gmcCC8zIZRP138fzQFaXHvqFJsN/ltE+cUrS2nJ2hw6T82OjyYWvaJsLbhjlyXgjrgGamEQlpRIB
6RvPtmhHhk1GOMbfUpDBCdsMDMnSjXlbYnKC2XyYxhCwk+azf/bmhaso/cUHzCeeol4szOifk7su
BWTX6i0s2xqcvN7Mud8qnCbjySiKDqGHL9Z3tQ5P+Zsjp+IRUQJAQP/EyqNWe+KHnsJvEVfTZQNl
LgA2yF+BCZuoJLOKupWTniSD+ScLCHbbwRWcdA/yAdlIkIw+ffB31dWFbDcVjiTkK0KU084ciYUN
qo1fem/+aLlPuE1IQTNdEi3JcXRWTo/cXuxNkgo5h7VL71xrZ583HX91PiEmqrZRcEHk9GaMzK0a
ROAGrUtDLF54rfsXty7CG93wy66fGAnfsn692XmJ891vrjImYLnOsLMk/Ihka6oR6BOjr1irnG8I
OEv1gYxzxcdVWku4UXUztA1FOjfa8kIFDhnpGo8cMZZrwxe60yoGmWihDweN7oGlQwrWBWoI5exu
3fp/PmB7dsmD5wwWSpFV4CiE08O/DRWbwaATKwqp5GWOu+AefZSqcMVoMTZf6RSzVGTtyOub+cKP
I1jLero533qqUFAsK7lHy3P8nCIdIdsmcNWcj+DhK3k8McZv5DUb3/SQlrYLLeBrZmINr0PcN6b/
cErmS/yqmzacqwKQ+aGs32AW3xHImIIVvQ0b+jRuA5rwtLmJTqEQ4EX06Scch38s+i8MsY/z4mGD
kUDa0avTEETanMe769Hral7rdbVMEMlz4AE4HdnYKrGecKFD7TutfHKxn9Qj9kqqiOHaNhYStHJ2
Ulvls46hVxJh4arzPes3MOFRbYKVtXOnZjrZFHkrla3TQ4N5R/XTffsrNEznFcX5WSSuJKzvD5eg
wiWPEvuYQB+Sl5NQdM7d8iyDz4P27cvEK66cmK8KXYGx3r+4IMddU67l8ON1wdngKTNLYd4iicyf
xZ2FwAfqyyWzIIqRLKZAsmRpXYAOvTdnLp7SuKJJcW0Gs76vphFcKdXPweYl7mjoG+zNMHhYnR35
xo88JXUCEx0vw5RckbXvgyH5+Tn0Ks2TQWFS2q7Il/afeXWAqdPF8S+xE9pppOXU7hYYPT+sI8zO
gaX46fIQiph1jQ1uxbm7WHsRwWrer9MeaI3xf0X2am3fgve5VuTpq9PfboZIz64ywGf/olDZbjpl
+fFyMVLHMQUG+tU8yK6sxY/V1+e5cAQ71ZeC3lhTlPTja3rDajazxhOBPak5qhFLY9DducmOf9Q3
Oa5ux+Uw93CrNS6rAjiK3t7zaxCyeyLvEiGwsL1WcLo52Tb7FVnUT7uJNmVtn1QuLPB8hiuc5pWw
VQG6kxKFP7Nz8iGCV1UcdExT7OkGNlWc2RDmAlcgAp+q61BM1Nx0zE92G0eyF6vNAkQgUPU9Lcll
eiufJmlpc5YIB5WBN3IghlZ55vGpZ0oRgauQW+yEicZcjrtVMb95hWhd4TuHxrx4N87HqWYwElmD
9OLkGO1uXvIzcbTPEHIWvWogJ6POJXudjm3zaHD4t34rPzJECS2RL38km9rb+1942ijf6+RPv5Pw
zFRUr5v57uAyKSnWE/Lo71tUN7Grl0ipvfiDjaiR+MForun2T/Aa9VFZS95fvOgK4ggvUrgYzsPH
XG2l8sHUZ2m34CeBDloR0E6OZXJj04W77SR1Lg7IeDYFEcDECRpch+piXGH5GrFopPK0ubdr2aBD
MTgvsrl7jPzWbckgiOWCKs2royeco3RMyPXWCjnkotR7q/3WdksnlxcDX1R+2lUoyKsRoFNttzwc
tEIKIueS3G4qMxDEpy+J0V8N/Mh1w27sv4CpnsimUeGwSkTkBP8DFuCgRAuVqeW9zFQQaZ3O/IQK
WYJ2uTnsUlCdjx4d3xC4jLqgdX2h6nfblQeX8RtoxdjdDwhcDUhdDoztGN34y3jHJVUx6j2T4Y8p
Sw8cs7vwM28xWrQhLyTQTobJMpidQtust6AudjSpjlHpJw+jjLuSHJJkIP1YPWbsXkaU8MUwEdlp
ucHB0rDD5l1SudZbTgdSsQuFzX6JdJE264V2DpoqDHkDjqUH1zo7p2sCeBuiid7tVknrKWe9a8Tj
tvj/n/SDDyAApVDpp+enUppeV/SHGRJcTP5qKo5UH4gQ5ZLLZygU+8nCmWWLiCfOxqfkuMi52aJ/
ADTr2HwrsYPcS5tT00L85xRATGA7fTmjYZfeJ6CDeYW2VS3LopX3RYsdrmjwk9RFJVIOzXCDqGmv
QoEDbUAyDGRymUn3D99+wETyy2M3s+zyHhwXLjtWPJqIyMLB9uw2kkvrog64h2mwJ4A4J99QbVVM
pHAPt0gVxx0iuvH0Wy6h19RiCjsmiMvUpvgKXcvz9H9uzv3NKLrTCbPENR+3huIFTjyznSUS6RVS
7kmSCDW+qhzfdmgXUwNchHEkB03AXAUSFf45FRp2V5KMDrjgAi97jdLwaZ/84AwPxSJctJ73NUtW
G+GryRMq+EBZp0fqiJjZc+JlgEZCVXrH58KhpavtmyJOghlqRexlHA6bZj/bVGlgFUGMXAFDYFis
iazLMYGISoAV2P5x+Hbx0nvp44ibzNbLggtGYJnhBl/uH/AZcf68fXbgAZN5dUkcjE3UA4C/AFP0
iV/z3fOugASghtG8dmct4JuEsrZDCXL/BlYZkMbctC5TRHW+dC0fotMzJjmFtbmO8NNwVwwiQF0i
3tFmfs+pdOxHLI3rbk4sxdjKYOx4S9cCRKoRVCPKG140TFtFnHDkn0SzCSs5ct9JmhN7Wgeim2WG
cTD0BgeeHqAAVVlwTtvqyAtn/34ySoohKuJUEOjCCCLQeNXY3XsXw/tZcWeN6mjuQE1tTMP9j9+p
5BZF6j/DCiI6hue5en5Uy1UqbjbqJLiWemo/KrSLrZ/Se2YU6UoHycch77cfRSZblCeN427q80iC
17Bb+2jAjfjooWACAGmPl2LNHAdPsOZsINfnd7sTeoFFBIRYmW4++MxqXHtc/Xg/fTCLljXT8HeK
n2fQr/3eFg6JhTJGG+5cktsnyBWPozW0inFEahn3r5VkF1c3j2I8DuSDBkE8KNzr6HIFRt/Jhebb
EmadSLmzzdAjdJGWW/0+nOrpQdoxiatO+FEtufq/CT5Sv3vRi5RMI2D5mkcbDmeiMQNQmYZuZaTl
ZyUNS7+/BYVUR8H3rzFqTKdhzMR9K2KA9GHSc6kIBI7YDDn0iucbK/v8RmptzOhOU1TJvmvTdyK2
9yQpN1jC/zYeGWJjn5jjopOZ067ODdrSXH+SrKv28L6iYIi2H4woY+9QRv/se//iILJkjAhUCiwF
a0V9DrK1IX6YnXRe0aDKtfCLnIenIfF2UOtyEX0yr9bglO7sZTKcIxlpJW4+QbSOZUqzfi4m+Ws8
u9W/OgtO9lRAjG76b/VspPV1nhYVLqsOBcNv9awwq30lhNY1Oc5ZrypHjhjnQkcGNZC27Ctome9J
+mQWNiYsnHQFtYpq6DwncqVqGHsxCgMonRtGSSHBbBKldYhZZsNSybG8W4QO/Qu9DmoO8hb3QyTw
ydzcXlaerrYB0uUjkVWxTWmBPs5TNzBnYmbNbGE/Dv9iu6Tv0ME35dO1Rl7I3Ln1E/YG3Pux5GH/
iHwWkvLVKmYlukwyaR6Eh9UjExCKAxpcXPBYfZDykKQZ3hiNQSaiLB/MRg1e1MorhrMFuPB/bCuu
PsxOLIGQXS3zxyt1NJNJNRvzhawokgHvC1L8iAxj+Zo2FMnR774VVnibNt/C6BvSSWnOdWv2N9ho
M/NP4tIJ3q1n+tw4TFK2ceBZnPPjN3mz0xfJFEoMF8NKMjtuwyufVsArYkW9DOeVUtZpjwAuuzj4
SYOpoAAD7CNfsw+sdSLIGy3Xbk13YnslfKVZxPXEovVkG5Jf9Wf2mdjzpvbLXFDkigZ4HzYtu4bl
nmUQ9lElzayVEcDxGqxJ2Qpa40K9kptUDRJN0Lz23aze8HO0MoaIydbBXH2l6MGWN54lOseBCBtI
4np4v7/p2d+LwvDbBm4lv3B6hEX/N5SraQ5pwLaCc3/SWOQUvczmg0cUaoUsSSXCyj9tzVxsROY/
Hf6ISn62DEW9guEWbIypC7kNBtMjTLUo4pmCGy3vxD2IF7ava85om/PyQqeV4G9MkscoFipXeEHS
EOQmqLz+5iGuoLFGLDXpRSOAJ4T3kPNvODeOAdoH3C9d7bkKocNHsXK3fksnr7vCvB9d8WMgjAsq
YnSudviWcZB9vpa2BGsDyodmcZSfB+kqQDYF/Vy3IFIrRDZlGe8FW/lLBsOa+nrrFuiAMwfTBDtl
fFVvUipsHDnXOeVqyCSQk/jqPS76BKdegYc45vnjBRsTbcV1GBsiXeG/4+ZZ85I84/AyBTW6+Hi0
r9WDltPJrTiDWOrfdsOyLHEchfS0ULKsVTRbcEU3XcCRV+0PqNv+O0BthmHMe/mNeBqNzaiFZ0NW
Ygw3sAsYdAqOdKOAJOqSicx0want0zYtHn8YYL8Qk3qMGqL35GbhARogA/VL6+DjfWtjN4K/iO6t
GJctsTn6hdaeRCyVNUk5GhrrrhouKVujECnUEJSku5iAI0c/oO7hUGExMx19ESLCxplR6Q4NBcDe
+4hxO5JrxH0ruznZoIdJi4BJM7CfHV3K+EBeKwBX2JtqP990oGTwm203W0wiWQ/ljIrLxY85eZrU
1NAuxqlz0TEsdvmswuefhOdqXYKb834mw7n3JC7H0rOyE3p0JpX3m9vvk4cizk0a+TRGq7eWnxxV
j67TFctubYl6Tio5CM9OA4J3A8gm5KbrU5EXZmKBGm9BtYSNB8UyCE8cvhs1w8OJpiUTR4PCGqvZ
/X/j55ZX9Nqx6zS3VI6sYf1oXQWVDbzf7r1GMMeyn5+zn95pH1mVG3M/ijyqHi63AkeM9Bh/Z1RL
NOTTe5gv61tk7EdISvjk8vn19MiUkETHON523TgXk6cVtdfs4xTSl4nsH8jc0b8YxypVaPB7erI3
/gI5GXA9Vm+8T1uEWOLu406f/prhULIrmMWiUf+tLHCq67ahtcKADRwnwzuLCVDI0iYZEJmchmCW
lgUesOrGGOmhe8j00D9wJeO15E4E6UdIrbfVr/WN/X6MukcoUiD2HNT48qD/afSPp/on7e+0fOzm
bogrcjQg925QUs+fZkgo0aHc0TzSNmPv9o9UlzeThHGF4mDVIBMxAlgj47jhhd0DAAPmIJ/t3Obo
d0/YLWelM8ZvJu5RFZcPpT4EdyP13vhT7nkqOtf4TDXL7rwi5N0Oqhh3GV6uguyiW2HOclzRgKLb
wNNUdlmFzOVUQ5wDFPia+bv2BdeNZzHhYCbML2J7poh5U/3WymLWHkmsw9nWv3on83lVgiZijV9m
/tZZn8CQUUC8MfjwWJhukSOYbReTRGI8sDuLhOCDoLRqYfko/g4zNRt8UD0QMkgqzza+rbneqJKN
EsYtwNO8HJnqd3Ls5Eq2BfjsrijuyDAoK1oYy5txQYUqL+aMJocpl4WyORqfqtJQzxlMFTVuurkf
f3/IXG07ypleBfr/JG2w9IrVQpt7dCGM4SM6aqX0PrkoRZkEFm+8cw0SvRrPRODHbvZ2MtL3sK1T
m/9kUU0SOnhLVKuhsiTB8QY7xMgghTgXfgUbXXcMCE1xHtdXlmcgNFwtSSnrlLI8MX3ZAZRwTM/B
FSEfSvGi4IajTcPcJGdZZWz+4KxK6yV3+udEuMJy3N7DDSQQRKaRfcRBmz1hvVImFqiekQevAqZF
wUQXX7gyw4FMogAbEX7YRmQpYc71ErqwVotntTRfnnrR8qnZbMzrgPPGLsbf7S1TUT9X4Ir3v+7W
hhA3YmEXEayp3aOMrxhF/dQO+1V4qrOA6ljac6eIr1duRv6B8rHfi21bTD/dA+Iav/yefq9C/pQ+
5f85gvql41390sLaxhSeQKlcW5WHGtxcoBS/6ibMCXRAcE7f5uHW5C9UJDOVmgS7mdrk1USiJm/Z
Tjmc5MBFe6UA9kzzKFzPaN5xmjMl68L0rXViL+4IHI/bUln9GQ83jNNBAu3Nzz9AKnI+EL876hJ2
yqZWRjaUDZv/ftkqfg+oLovDMBzhIyspQdbn3qZqYMjbRShmrFDC45qQ0iSSZx5ydG59Idvlp9MV
2HJ/g5sUeKG87oHDctY6yU5Ab4AoHAxefKhE3ZMK1WQbRI202WWM/5OxStYXMi0CrBxp2vkGss+o
p4MO8JbbqnU4K7I1+gw8uZH+T6+YCAZCT0jm+x4erukW2EFanORhtZFuFq5cbKKF4ZJAmNwVu5OT
Qm0l8ogp7DBp6VNiY4+RxF2mziSGzGHBlpglASbK1n9QcRqB1YuvctCWROFT5CWKipbJzPzpwUsg
0jo7vASV0f40MufhNgPggpkMaRzJDZ503WfGA1sRdkA71GkwnxEbxNEi/OAKebkQ56bAqKtLjwpa
DtgPBFS37fom9/6Aime+k7pw9ZL6sjd8Y3U1R8PL19FJwtr+H1F0UvNk1/ilsT5htkBWhooNQnuP
87qwawMWA118kilMZZrDGolUhjuaR+CgXJiQA1S/ky8Vm6xY6PKD68/Tx8UHqqFcNaadmBG80x96
i6OazfKwKQBqeAJrTRR4ugrUiD3oEO9Ye00+U27F6AOheHEcQ9tjYvkJGyfkhbZREKoErOT12c8a
TEuzaxO1fWvRjFanPjZEqacPWSnEzg2HC74RcfOZWXzz9N5ZRvodW7H9VEXGF2jF41kfaCFeqJUB
KGyQfy/UpUB5ZcgOi5xBMrfj62kgj4FJTiCE/7kKWPA9RkQdlPf3yBdw3Qt/TnIXjRDZc4aPSK2X
HCzpXw38aDVnMO+LjFT8un4iZuWqU0xabHK5F1eHhAOJn5KpDPKtbSLnbUmdWmDSSBgVDv2w/6c5
DIFBBRkB8Qr9S+vZmTcvQU3c9G8SMj+MsFXyt9glPEldpwAapqTtGSEULgd+TyhCAexN41UqVKzj
4zBuSFTd18ke9zLh8JVjEQjzm66F6ZuUswtXtuYwSgzqb0g/NM/H7iUZqfHHvIsnSPBYH9XP6b63
aV/YnpjYve8tb1ULTJ+Xlb8GYjTw5P2Yekoo6TtAijBltPRUnmi9DS75af6F5raCW3URlD2gycsL
UqP0QBXJkvD3Z7+9MrNymTKqhEJg4unp7WrLm54P0dM0qCONvbpnHDSvFD4SE08DLRzF2/TNFBap
0g8iSnp86YMYMfuLErBw87EPC64xmXE1gK5jkqhMJBUKojVxvi2syrFSRryhAD5ptTns9OAv8ya5
E9cV7k+uW+aYh/FxLI2+3pQKUzi2KyVIIQfmRXPZD2wXAExdHyYrTNypDwsaAF1SxiP4tC6BVRBX
41CnSrpokBf54klPNjcfs77l62cEuzakSaeD3tCxgW9+bIlGZZ2uQ+uzBW4nX0+Ur399MuDPPJNf
ZpnUhjqiQQnRPlo4QaZpswqrkayYDyfjMFkbMF9VDmnRv3xlRaW8a5vGT4n70HTJxXAoNvX2bLak
4ZALHayZqCStwUGgylrVRTT1JbeZ2DU/UWBZqasnPvRc1nVAM1C0yECJhvRODSC1C8oDlX/jBql/
48jtgbenLhq5V72j8FbxkPqzoXzG1lnO8wjGvCypo0Ve5JgghW9Lg8FpRjUf/cDDfSv8kx9ruDtR
CCTnTVy3muAyZYkymz80/GfwTiMRElBY4Wg9m18OevmqQBzJHj38/A0ZsmU3wv5EsIc025OLRCNc
M/JnJQVCpRYxNT32xTiBbWbvsB3lUWfgBxGuGvWB2kpowN10np68O5Ji8cJ45R4DHtjIwt936cLZ
Uz2+toNPVbvQRJkEjJwfmdLv6Jpxp7nPxGtLN6Xcon9M2ceU63Pm3ermvIz88NkWkAqafKxzhDdp
7eJZ8AEdmPg63BeNbLQ7pdv8vPPid8Pkz4CHMwnkFh2nU+AW/y+qgUHQMumgYFV4DxMnON8ls0oH
Cr5yJwXY4uECGD+pmQGtEZI25WOLY1Vf6vGLesvrs79tlRJQ3mWq95dyiUzPyJenm4KUyDWaYv1g
mEKqyYdKrrfytoqHEiP82fO+osIWUQobZ62RP9RuvGccHQTJa3/VIg/Am7TC0eCUpFaRjm09Zet5
tEo9KKabjA7n75QzhiwtKSraAdjusWxvp7tdftqeEUH/fjIDJrEj60mJEsK499KbRB8tiRtkLEwR
ItTTfCCS6VN5yjeN4gKGkbLPTYYq8P58PMmwlC5PLwXGIbrAz26wbYVVgF0OOHzRlRHafuGU0kKu
l4owhWYo5/XDRuYtkU22OHRddXwYzUmrohCspjbgKxIvMdxGoKQ0QFWMbyxce/eDWvVz9555mrxj
N7Dn633I2XsjnGzBhEL3PeThhpmnfUBOvXCtTHZGUMODw4eP7GMpex/wwVuOGnzisEPFvD0Lflbv
L5f0pd+sE6+KoRnRVmvRJVSBGBCZYbWr8GbFwsSUss0wfg7HU+vBDXX3+OHAb/We1CTfLSlf0PrV
i54rgJVyUHP3b2wCvfJeUu5O0bXDLLwzS6fQF0yoEDfItc8h1KoZ7tPfD561VFkFxUG+26Hb2wI4
zvLaW43VXqZJqejv2WzqUtBWTvXA7nFDKNf+kVQeVMEO4BckNIF6rHGOEeOlgQk+0E+Q6GLEBhvS
MgtmuiY41dlxQUE5lE0xafy3NjksPeJSO+qgeT4ln8vAEKPcK6oQ2Bgi0vNAlKX17Wk0NmK8UFNH
e3aD6Za94mKtlW8I4Fz5ctskNtKxRpuO7SZmN/sZjSqX4ZMAzQTZY/mkIJ/1wPaJn9kmicVo+JtO
DrnVA/ZwJttCN5Ao2IClwvEKxDREhSy7pTS9Z+jmbEsmAdhLGr+xCDJFHZSlIsiAA9K1CmfkDz6A
Dy+98FA2LwwvilcNNWYdC8MlVCEHTHkTrRxBRtF54nGbxYKQmNJFAqahPOBh65TAb0+X9QPeBgPl
wE5q4MPwScDHQr+J1s9avbeL5BJDIvYIkj3GfeJgINBgQk3gnUoOYfE7K3/0sfIZ0aH8rIWfM8W+
pAGnwQlWAko9zB7841BDwvBu0bBkJw4pRdHns5b9zIOnNF2he+fYGIba1zxT6sHfXrGPouSv23Pz
2VZ7JnUExM9MJjho7UC6OAxf2wzyfunmH/QnRTpzUCw44SzHKOoyUUmRXkEuXhNilcmCxJctC2D9
CH02ANgv5E203O8dOH4XnWzihB1O7lE3vBo6xDrd04mqrFBvb/U2uWIPO2dWuYusuVpBfcpkc5uU
r3gn4Wq/RcLLmEGG1gI4XSpitXXPUIQ6UFhuqQWJjf4W155hKHfy/ElCj6kKcBCsyzyf557nJ6Ni
vr0fn6ek8+WcijqgzklOttGDhGFC7/rw9n2KfMv4f1bm55vWErpM2nYsrWaIQQnmGtGKvW9MVOcH
EnZIUnQNAumHk1AXd+Bq3aNlzXFvIwU58SGhfbnIby36z4esczSa8m9nEZ5y6LVqHGxHl4BBzQCu
0wKKAZDAwrEpNdI6hDPnn/2dxLkPE3pISLAKfHbNE+bJELUvCKOMXGrDPp5Vr+8II4hxmGObG7Cn
UuXnrRi09x/ZSUVFhucRbdr7CJ/Xe2KvqSdS9b69g3TytPiKdhlc268bq7KlCrny6OweBrK76FUV
Y0krVRDzhZPsvy3oXanHkvF7b3NIyr+Ntwzqcle0Ur/JF+FCXEBi+bU4GRMphviJiqm7v3zg/TdJ
kGxRf3IjFCqA/FH1JidUYcd9Z9KFhtC/mAE1ETir91xIn1AHx/T0FuD6L3Hx5erqfPHy23ctMaPF
NOR4uA3i4dWf4JxmuxsoRd0kmPvOJmnaaQVmGBugyqGIrPrh86UMB3NnVlDtx1HX7CGeBK2aU8ng
bjjfmFHTXW0QOkGruik50M9IDCzsr6DcQyS5m5gypr6fJgOk4n819hyfERutKxmCm2bTKPYWcehg
qvCEzFakdl0gGW6d0Go4cFbhos4SFofAv/FGdN/BZXFnI2/HWX7N94Vm5a3xB4kHLB7qeoli3Cx3
o+71eFbwlCshBPDF17g5iZEOxu56ymseRFqn35qIiHjbBqrl4hOo8VUp4Q3rrl45trYwOEt9mMGH
hqO2pAjAqniTfisn+G75g0eVMGTehVH0KkCUyGzHXQWWCCXij1JVck7IEAmEPvR/2kF20V72U0fx
pJKKqR5ytV1bccTNuvS1yG4Mbvb73nyMWAIkXifuB0TD1GGN/b9EOFT+kAnKF8Dl2x0q+YIoRb5r
DXwb4jZ66DLQ7Q+4FqrRj/JK/35c5fskh1Z1YOf7YJfwQVYJrAFy46dUCeJa/BWq+hAzF0QJ+gSk
cFaub6AhsWANILvUHCyUKfWw47ggYFGMy3/ESrBEB9Q1j0fplUkBtMCLyGy6xl3ubiYt3F1/FGgo
9gy0wQBXb5FEOGH9himxopFPWocYdq9lDpa1T7E4hF6jQ2WRqDsZHOqLAB4pvdhovkS9oOzYkUy5
/OXjX6dOJphmHWTosrrrkRco/iTH6uTDqx70mDJLdyhb84/QtG3t0YVaICDHAdrdh7OKGKDO3Wvx
ayCY0z8vkcQiONbhHNxyKKmIYqvt9oSZjBtg+8/UOOl6IfwFC89KHv9ojZ2gvydeILHjQAkZPERx
AWSVlxonGi+IgnUsC5WinCy5pjiOFSK4GnWA83poav1P2mg/44JHAiRBwXQjAUVv3008pfaDoVrL
kC0ZWgqIBOrPUNNAhLDjulJB+GHpMNuCNmYoT+ZTAn7ta5iTl+DNOPq81OnovzAHi/+7bbrFI0Q+
1TFRCbQ6H2gBcDWfnLsulvXvOMdAN0zcdrsXkPPZ81Vo5jA/k49sojD2nPk0tiYHIC8lPrn1iw8X
cwlIYhw9qnCCaW9QCr+w3rQ1FWPVfleBBKXxbgzXXSkQ/8wWXNhVAi3piv8YQs/F5QV6V9H/c7w+
qtqv8bmDP4p7NKR9/siWdCPQShF1UJqWYxYWcu73qDph/kLcrywzlvT16K5U40SziG+MuKxNndY2
U2LADAop9HB73HdnGziLApee6LvA7rQdwUhb6PLebhun6M1R3bS3bsfAQjzLJWxuda1seWxOFyrw
XicRn+YoaelaEkFbg6SUk2n/F44Xs/LzA7Qkj0DCgfTiGDkL+y30ddHIeIxGS0r3Gqa0sa6oDZfe
a0YynCRbMdXeVPgncj/et3F2zSkgcb7GSg/IutDgcXN1zaw3aOVQtYy+wUGVVV04mCiMYyFQHwvR
+FDpRTiTqHVVwH8sf1LQ5d8UBlxl4dVW4PhttoY9SB/T4I6nrw6xVlQriykokNnKew+eUtawyYPv
X+xOFsKvXQBdgwnjjq4W9E7ZyEFRVFgzZ4zMhiamQeYKDfXR5m0JiCRjDiPspftCISj8zS4TZJ3A
CJ59AU2AmhvMEzKEUSxRoeGwG0wmH4n3As+LAfQEqOfb9/xxvZf9CwrFdbmZZtqHw/GHqBFlajC8
dmxfp6MWF75uQntWYYuMBXjZsXqUoWR4zGqSPePk5OD+mdno47jwPBjjOz6IDGieEASCZvWGY2e5
N/KZNPN5C0qwQGkCze3gCrn+nFs8W6zW3DY52kgrmPJpxv5E2BVDpUmZvr62CdfRrGlIPW60zDCj
pYP2rR4RfRjn2mA/HHpZRVsAnqoY3w5ULxCoggx0dPqR8DyiSX5JQIn4qhOPsAFSYuYNhs1o3kcM
Ylhtz21gQg2aJq1gukFW+rT8lyW5vYCe0UCIqVs9y3M3U8NR12rTgzX4iZHV5WCgvKhYzKzTakkZ
HHZP07bcCGU+28iKFauOZUeDEoemlTA23BX2LPLFPtVgyS1STz+Ywtb8OWOfUEIM4b++SY/cEcUu
POFF65nb+v/qa7++CA01U2AJl41KcEK2E67tV9kFHXGjaBzJxNKPQIiIlO3u/AaPsH0j91On0q/E
791yTZBFkIs8N5Fc0UNr7zU+crz/ztu2W9fxmLiqPRfcKZ7fivbUqMgHr6dGebgWCLL/2eQLMiiU
tmLBuOBkYZkS6UhVrTwUC28pkNu9rZHJ680ab2DdTilcP0XWbI7S5OkYZWGTvXPqnxbYXG5KgeZk
3j06YoHhaqZlpbSuyUxjGjqHbZ37d3lh3rSw+sKaqS8QFtqgKyAv5oHS/NqEEznNaGgMYT2fjtiT
/NnFeOUNRdrTfAGd82f+yvrjT6UfgZQAK4SJR2z51K+HvpOKXSVl/FgTe0ePt0mn77aC+JXBqw2R
z2p4gmleuTJzt2nab8vu2S5hHXt3jDoPfuyRAtXdoKEtWH+n1n33B/g4HpEsqtgHO9B165f84yo/
n1/wgUNUZJiH/6fjS7bY1XouLZtTkn9uW1gbdyx0XXWjfoGMfmCAU1p0wwDxilhWLeclSID62Y/S
cJLPmXpRsWq1tSsMUxYxzux/UweAF1hQq1yhno5dyQ+K1OYYE2q/ucA/DlNDbQjMSGBVOHls+ZwC
HXfaEYJTIQ20PfDEwN2iaoLg44ED1rx3gL/ZJVmU9n0+2xUhGqHywhN8as6fl8V51UXyFEJFBKEz
rulOnvVM5Egsf0pXwcHnwNluA3XFPGYmV0iV4ETGbJLgNPOK5dZGi8rQ9NzED6XLqRO5irO/otvq
im9vtRpDTpwSxmmbJOlqsRxRuTHOgaGxDzyQlhiEYsWTSiyp6aSLMu+OK/dCYH6aONCu1vhcRPmT
L6kE+Vo7gEtueb133cVEbqgCVqSv4nwwOSYLrdVWIn2wASz6Lflv1w9/3yHox0YNQNoPm3v5kMpY
SL0Yz6ElvjPUGKBFI+RPRgbsA/rf9QFTHsIgRK9NoNeeUuYw+m6U4fmGQXs6PFMD8FAED+YYo89K
a6sB2Gbb36535Vxn4IvL4VmC5MH4VM7nozomqWDvoMy6chCOXVpPrLOYCDUi6/00lhxb3R1H0eUq
e242TozBYra1yZpMuHYGj8bHaBF668tZHHezPC/mK+AR8+MXZWOTmprtkGK5nA6GTRl4K/LT1i4h
3pMFHk3J8HyAljbyYIvym4Q96VlHFodMxaclYJNWfz9pacPnssvyfrKAQFaxb9e9kcTD4Ct4M4gJ
muwtkJA4Rh3f8Jdg9IdkURbDyzoEhdX8+8l+9WxgSzPHayUIWfv1Rzw9/iZoF++s4eL4717uXKHS
CQd5V81K5EDZWsUGR0TJBIIgZXv4V1Imhn7j79lxWRpOPhsk/stqWiDtRzClDZaYI8m61PNNXoO9
4S9h+OYip0AApFrKrAZ5Aeb+/Hphbx1VJMR451KqZHxK7i9xiareiV19v5wDLJ+bkQpbWclbbpHQ
LvPF54kpKeSE7IYNhb3xbfOZrItup60gE4xywu0qxwkGaMRevs1fKJMRUu+EHAG3sbbbOSi2+yzJ
j4ViPVzfGpQiK0d+agC+1bDE9/N+Q9EhkdiT1xaC48I3pt7f+NqQqy3vW1ISNyxu+RWTQRw+hweU
XqaHrDjsGaVf7VrwaolCB+HiVAURT3lIErpigFR5t2gMImCWOM0Z+hVSY/YYfB8OQ7jzRen0UChq
zWLwOiaSijdUxO8xUcubxP5NTYzCtyy+xqRacr66CrH+AmHDl5JnzWqT86wOyLcd/R3XzoPv3RNN
+EW+LZWQ0Bc/c3APb7n/qvMjxDChkyLZ7xr0gKr9QZZOtTgT9IbWE3d4Rc05b5W78Vn1kRLi0tjn
TkJ5d8Avgn9BXcaysPmMazh53/WPJPB4HPb4YtZ3sAaVTgJEGQ1emmYx60qJf5cMFnlyBBGCmHgR
aGADms9Qg9gRDv4hZu08Y9SlbNMaJigWzH31JNnpVPSDBkZAVwbWTc/ikdaefTvNCXLX/Kdhr8L5
zvKDAEQH4valQLUhT03pPra/+nXJ+RgLXNgZ1CZ3krgNVD+jCVRDtfBODSQxuqkdsV03y5cu6zdU
Ls/ZkqKoW9DFnHR/dXnMKYiZy2XBAbkdZ1EU/AboTXmHHBMJNAq3D9zpFZalmRWTU7ueWYAgOe14
TDAZW7z+qfHh71ud3+C4W1HgMMF/gOOdjCa2nR1QONB1/SB/9HIHXHXFd3kvI0573a9IBMW1yLbq
CWpm0aAS928xQG3PvO4TrVlgDhEqFnK/NAiu4319dn7nqru1vArtJK+yQOuDotzKuN/x45BxkFa4
B22fHY8bw92JVda5wn++8j+t6A95hkPaBr+2jYuctyFWtcHULaD2AUDMGH4RHXulFKoPTWhId4tD
YqCARqy7dzBLa1I0qR2QEv1oAnuwY8i6/F+dwEaH6xpSBFFMC0TE7eCljYGvjrujqYKD9isvI+4f
YghxJHyKVWeH8iAxItMkfqUmRyVp9l77VgvBYm+tfchN1jjGr05W7MHMRpEF+vcls6wURCH6FT3E
53QbwDpSQFCgR+nOUWvQZ3auHHmU+7VClaWbS06BLrXzWfgFRSjGjqbdG1iNIrFp5ccb/kKsk+Y+
skv6myAkD3nfgaIpoa/+74clSFdcWyNEf76MMeWz2UEJu7qQT5EiMRxEvK6kLAlvKMWfgQ00Y58x
y8AVyIV63Hu5lxVE/Fh3b/pFib7s6RG0CIw2pqoRC4+NkGoiJ+HvIzNIi0v7U6RzG0p5kuW4P3M/
jrnrAivrMGT6210CFVQxGTZRCN6Jgf1stU2LCxaLBm/mnebn3S86du/mbSHAWOivjKVk3Mo0Ou6/
KmSJvP6SY68lAXBU//SuUuy52wmAjvdXuU95MXar38nb4BlPmUjTXkM6iL9n4D43HopdG+y/CZXK
njS9GjUJf7h7pARX6d90fTVoAuF4hUGEDMaeAJwxGgUKuDxEt2KUbusX3H5Ktac5O+F18aXt5Asx
CNM36Hm4ltboAWfXnTI8i5/UaL8EZDFjJU6EgpwD6b4grVbXgNr7Q6QrbUQQZHSYnTrPYy2HN+wA
xJi9wfOrJhzDAlQsXs8G2CNl39F0q10vJDVGkFLjBOp9dDp1vOsFJjxy+Dy5tfTi4SNzSSxksSAC
pQoX+eZcSZ3oimSsLspKvsrK9ZIdIlUbng8t86xjnw3Gkp3uxwzZ+tVFU18RFb77fjjIHSZyteWM
LmTlaU2XvitFLNygx5he+Gbgby3vJtjUI0jA9R8+/uQ6JguU8NQgalICsOR37r6dhuIU0ZXVJPVN
F3RLUsnnR0B1IgTLEJ7cfFX3w1dnpInpzeDEUOME8iujS7/pbQiWE9O8RzpfsKDRPlZKZRnWUIvm
QYP4DwU=
`pragma protect end_protected

