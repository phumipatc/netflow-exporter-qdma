`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Um0drLTXPFuLHI80C5s58ILfkUPWnFif/3xG0/yjnQtDpYJton93Tk8LFd6tRhSs4INhxk3S0xQe
+TIyE51RjAbx6LTRa/moAhHTlq+bmSg7KRQtmlnQGota8BRaIivSjGApTJD/sxf1ATwnYvHK9p6/
LNFPozBKW0x0pi9MYD38aj1QzLsiQklFFV+3bISLLFbz7WUTKMAVw/e0fIY6zJytam4Sp7T17u9G
pdACpk8CIjpBv+7Po0x9CtPQBfxF9WOqH2rf/mAju8NTlnnn/ftgoWdEuWn77S5ITjv0CXCadFxb
+4ZZbsYOLs13P6R4VJckvBX201inyxIBWxkE4A==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
vYQzVF1SJl0/2SQBDw37BeFlqjruGDqFhVvuGhqp5Fwy0rJRVsFd/E7ldch5GstlrEccFLdXarE4
M5KulUVwQ4I5RJcV0jmXV+gRfphqB4p/s/DPEcw4kcpf/wJxDIba3rM/PQqCevKiyap6E437Rpp1
lOLPVyUDiY4kf8QA+KALM2jA3w+3qZAWsThn60c+Lim1BrMkz+NpJPzHI7hi4bUgwg/jvgcYzLdl
xVPze2GThmR+HTej638H3AYA0pFp6TIu8DeiDHFntokoD6IbhmKkLMlgdkeb8jixwGevGUiLX4pn
9bSCKb6gMOsgAp1O4IXPyeqnEz5qQhZNZyeSOgAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
nvWsri7HFoKC/D8HpzJ9F06V2vPaRTBaklgOoFe1Q1jj8ZjDWcEKwdVjWuthd7mp42eQdtsTTC/7
R4Qow31Ebw==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hYd3Z5F71fatbzARUL7MaANiKWLmfuvBDxakrUjkIPGBX15VbXnMy9dzOaeJDZrEOsepWDk1kqkM
sXTlRhXbhkH1HRYQjwyApXQZoyok6FLBYt9Kr7PupwP84JyATILrf7fj83BVPLUVP2mrGxBSz7km
dm6cSr8tIvQK3dh5UVAuJbHyEAUlXCK2z/R6UZwC9nczD+Amgh3ungSgbqMh/kTeEToY28v5BJyr
JnpTVeH/Hp0UeJcnRLq2vN2vd7AHMhjldC7d6apzzTv5Ifii1ZeN7WzQUhsFpDPBZzNFsq1QZJv7
fKuwnR4kr+xP8Xozcbez/FVRnRBZ45Q0hBVmjQ==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VVHbfea5SDOksGskN8Pg+BLXz/Hf0Sl2A+9cgmqHFAxXWs4qW3KOkPwdrQBqEGLBzgEiOMUqB3Qy
BYfAEShV/DNNF9LygE2e/IGD4RYg98DPSjV8pDYjUggbkGL9XXyZ23d9AZihCOZ7KBXeBYcWhq32
+UK/LNDzKohrYzd4NPfWOpREq7F8/H91usqJgwFwD8gsbyMzrA7LYMx0lSdC0JBbW4p6K4DiYAP9
zAP7Do/6jVWkEx3yr8A2jMX5IVE3XiOoVhs52cpiTIYqLaDu0i9icV5trmYzxz+5uzT0pVCq+tan
EZW2JsfjEmfuX7gL8Gq+GfbkH9SoI5w1PDTEyg==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
HONo282cEXZfvHvhWnDUy8ZJUGLvvbytZsgQyIksGr+kuw3zQIuPWtnpIxkiMP9fg8dDX/E1eLHd
2BvVUTlE3MNswiTcWIXsDPJaaeskcd4ThpEL71XpDaspcPz/vcrH15g54ZFt2xB539zoPOZE/snt
Fk58yKjdO5iDkfO+lBg=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
j4q6ypAQfFqWUO9fDnFlQCczkstejBP4WcHVDvCo40x1GpF+Ws1np702KfBfYTIcBtR5MUvz4610
1GBqiB5BzLLk+4c1QNj+FNEL4f5JwzV/SwFnWraOyj0XdXdibltnIrDEIxJf4CbLb9okiyew44RI
lWwH/NEJuvxJmGOLM7m264ugn+xI7dtObjevSt2GGp4kLCyk9v2tZLLTbbwPQK45NbaMW3Kdkv/u
SYDABe6my6O+gudLrZijlJzf+Ps3uXc9R7JEDUpGsmX8Tbo5nzlvIbMVIrspfw8WEqsb0pEL8U6/
ERNV6wjn6Cwdv9051/1G42x+0yVqhnD4SNX8xQ==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ogvw021k6S/FnwtUpYdYo9Out1Xh3iF+8gMm1vl3r0jZ8RywaqRy4055eOBhmxZYuxA9IfPGMOp2
az4QWhhev78t7IKJa5xW3f4a5K/Po2qYE2WI3txZSjB+hvwaUJKV31p/7Qta2lDnel8zEnkt0Feu
BxB0nX1aHZgQVFInptkiwIRPWCxworU2ak59mcSk9Oe0HpS//Yledfll2BxmJSnymLZot+n7vqxI
uuAIuFDOTLZ1XW13f9Ck9IDsq2j8wN7j8xszeOCWJoPyXC+VFIGjdZVJJBvLco/JEMk3Z6V4Igjf
GFfOVjukVDcyBO2mEbYawY56+eTNcYOPUYZw0A==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
MoJVu/f5vfn/7dXgZw8CoEB3sr47FB2vXGUk/CkBTXWeN09CfirrjhTGxY19ZWcDBipMKYUELeGS
9Z+NkdgdxTzg4keHcNy/9uPdMPn32EV9XJQZUbhpDmcgmDUW/ebRraLFjDA/j0GDKfpPJHv4L+6b
XrzTCuVc9wxHQRhEL5o=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ASIFbAM4ApS9iyQGXMED/cNnZQwuwdTrmjHNhq9B83bh/tMt47C8jGSsSZDqmY3KiR34xMofV/k8
9h64F4zkZc1hR0/MpOmfU/VyAzej0vaQ0NEdVkBhfb28XYU6A0XVsnIzJUeURyJFplcIL3rSdVE3
2mfCgMyt1wH3DB/IziL8sf8ovHqYikoS6aUmLSmIizC/qRynf3SrBUrAHmmXY4RAZ3gSOnEkXZiZ
A683fVpR4ariYBd2uJ8Ayu8IGFFYcYhlJArlH+p9Jm2GxVEY4f3DxN5GZvoESvslnWMvAXiW73Iw
uHg3YtQMgRGHi2J4lQfWL3o0FstJ5UcdrBNr+A==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20144)
`pragma protect data_block
9fNB6/4PDw5VVe2fJVtm+I2rE+ETPuusOuijh7KIK5MQ2RPdR+qOLa4Zw+9Sk3/8FMyezD0CNzMg
B3Z5RJARWpvLTfme+sa86OXfa4AJaUaki6iLFc/2S98FZ4qBp6yW0498dq0VKf1wiPzlX2+aBxu8
pDU1omJ+iKJCmKpiuiwduHy94QSIasq2JeAwW7HfC/SEcvSrJCf2lydVeCLfILHJd5TnFD+7UId+
hBHWretSmrpBwxBRynghKpv2XYtMZeBKuyieOwvYBEbAB/QxF2WlkvElCT4lwXhWNxmtoDIPLpT/
NTbTmz8v2lHuuN673HxPG0N3+eKEuM28AqWoXGL7gPZ4bxhfbVfHGCtbnFk1eivZr3gJ3Sa7BoK8
tLdt4MJg3T7Og16Lc6LA6vR2vPgs5WIAQdNpBfAIae4XbIxJGNIYhcGmBLfGPnoNc61TWDYAPSkp
NxsSh0g/nkQ3whHbSQtiziaciNZjHwPuYzDotNjT+dOOPaSe1S3RVSO5ctawsJRT9gDgcaboYusR
UNSGJ7HJggy11YaM0kL+Q3XAqAap/7wGxz+bOsxSRWU+RiCea/7pdLoS07bIjTrZ92Mpf/rnmCgU
+byVFQtCSztVXgo1E5/ycOASey3LrsFZeMCr7d4U9vQNax6aFST+bykw34jNocLrrp4Zy9TTD9qg
zMM0QPxq5QGjI1QXLvF5zfN3HaC5uqTU6dgv9ad5STT6ahELtAAm457lmZTlUMWVOWD6I2G524l5
EAoRrZWOubM5BHR7QdA4lj566Cua/a1yb5hv/1hJDsIPStQNNnbRHlT8XiJjp6sipH6BXDS2rJ71
uTUjdz4hBBQZKX4gSEnyWBE4+Z55IoQrDPruAKgmZvk9uGO7mZgzvh6DR81qM4ZnjjIm2HKKgk2A
qWjXkIfLOk7ziKMXFH4eVtlC7s/R+RzGvxP1n6swgNBXn7I1hj2EXYF0OhUbf5b4kf5J/0CVpWH5
aDix86la1dS5VRwuNZw4t+GXvK46XsU3DKKqbfrhKSZpSTrbI6bhuD6CVHzZxUt0mClKCISSncSW
sx6tN46yAlcjgBC7xOjHyMm40tOIr5WBbCLwROcbajJtrGqE7RolCAe9tNw5zbsnRYqiYF4xQKSp
wLJthqOJ4HerRHVsKjjZ7i69ltfmVkN/xsCARZ54u+b6wzc1KDYkGJXDFE7ArBCY8ibXRqauccQp
WT9RLghDMTsGq+WrwUpKxY85aSnKzxOQ9Z4bz9NsrIdMqxC9r9uLt9uqVUuYSzOd3gw2iJRWW9nR
fKALbt81uNgZW/FwkEFz6oEIWWHTCSS4uks2hqOKMn63FNb2pF5b7LWJf/KChBxTnJMFjZiL9KT0
3zVkrNGHck8AnP5jCF0RWcuJzOmxoI+bBKnepw2CNXRTkgSCBvGeB4W1ve0vnxKfmSoHvn7UIlgZ
C86NeZVgq9FLigsQGWGB27GQQK2iRq5sNxlouOyl+9000sTLYiky1M+fGjHuuRAcZPDBnXiAKu4j
LhfXGZWlv5c16GTwJqoIqxGrXfe8dG+6GLx4U5OjLcITWmyqfWPAdCsjzCujSyC7l2Yee7zqBrqE
0GVi6F8DHPHnfjBzAebjr1M1PrWldTMMZBzNKUoQOGM2btd/GSrQ1k8cTvN8DJpee4kJ+1Nw9qBS
SswAr/r+0+LrauREd2VhjmgiQuKqeSw3le9bIAlBhpc5aoy5SX9Mq+hemZ3x3Vl6DmEB4fBU23S6
jdaSvICR+MrAhGIaEc8xDKkG5feZrWzFmgueuKCqzGjRzBWkP+oGePwVTjAfSb4/FIH4WMG3nrT1
0aJaIeDwmhOMqsdNyiJo7qGawO6XG7DvhmErxAiWY8mV4vbZ7QvOOshdlGR+6FPAf96xcBgT6uga
04rdzjXIjLFcHgZ33ny5yxTNdSqgPwr+wjw/RjOEEmQvLJocf+3uTiTANhVTHKtM73YEQK8SNOnx
zXkey3vykz911ktWAAEJhAry97GMU3lWhwIt2K1+eUWaHeBgg+NhmtvFYuPWY+2vfJgfWjvXkif9
x9+ib5Di1Fi398afaOo9JHHvgoOr0NQYXxYv1Wg4ywmRNC1MCVaBU0liUjtZ3KfVazDiNamkZ068
7VmwIoK33Xsw4phPhkgAj45OYCV/bn8V8QyEFwvpl5gWiBlaL/kBa+edAKwoQctXgq2DAni3Wwz1
2xktiUx8Fx30enJ7G/+X/iCkDtYFnaKTyCIAXruxJn4i3TVSL00RR1l12DF09B6Q8mozYcRyO94W
DE8TH3HYv1x6RqbI7Y1ob6B9KOPett7OPxgdvtC8O09f7z6brOkQ0apqTrfPIODuBlqf6SziJZ6v
kIXlg+ZsarfKk6JL5o2X+azsoHPGlcpwkfWeecWQaf7Ufr8j3bhcraYJsJhPP4tgAMLFvKAssSeJ
NvRnTfRaNosvNWVnyReztCPAtsULviCv8ZFRmUTwp437H30IN4O0rJeUrAMTppQpwISy8LbGnoJ9
cuxzwOSd6dEAEurQpIcUFwXEwDsuHZbIHEsKxN/u2LilnIpVIzvZ3kLDt1HjYIeM7mq/3LJlXKTp
OtnGko+BAXuHdR0yAeY1SD/OujhlYp5hxjzNHoqk1dF6cIgylj53URiA8Wu89FmcGsXVOS/k+VFD
Dvf5pMhuI6Yz02vNF5AyQL0tQK4OLjie+RNcL6g/RNUFnz5Rn7muaTSJIhIcsJWyYWgmSy34MRjf
TH4AIp4SgfVmtGuvmt13yEbv6eDckmpHWd6Z/HlQPP1Hxr0vdCkgmzG4YwxqR4LY820UXK0QnH1M
1H4iMuEIPi0HgtgaoivChTSCYnwP0sjLJYv3UTv0FRFGI3hwmew033tDXkvhSc8KnWdHWcgB6O3x
9QmvHCaiVqiBjEDz3xVdEE9GrVi1vb9CVPVcyJYrVd/tR8Fj3uwo4N86GVu12jvByy/+SesKTsCR
ZsOn7SKXWUxR8WVgpRFSlV+Ng8R2DCTPGShWMPANDToKzf0TvlUeygLlUbVPk4g92BDvSlLDNUDM
QgS+ZJy3+1W9avtA/0vM02QLJayrlWV/tcjhXoFjmTcgTrWo+WgQMqlYZBzMCUf6GrJ0bG6oX5jU
9MD4Q9YltyOZvqAVyWs/9xcgt7jqWgLDfy6wBcNa7cS6Wt3Sg4GVvhg/BCR9CW9IkTmeE8/QWdNy
vK+ZWgnymm8iZFK+eL28FZ/z0LiAF/aNVmyg8z5vhhuE4VeEm6hvErhky8YXUzyEP8Y2SWGFp5Nr
z+9Yaa8fCp6vPxSrL6uxBocqVE+Td4l3E3FgKJJFFLfhO71mTF3vTi3uq8k0EIvEeZsFVrMHgWHj
7XYBXXxpcP9oUqvNgXUj381tcqmXuBGpo7EmEBpMIBa9sPpAjAB9aDyQ6l+536Zj/urVlOdQoksC
rccvNmJkLqthpRpSIedTWDP41SH+uyICh0zUuzv64t2/Rb5/EPR1M4wJl44OmtemboM3ht2oUhll
yX6NTXTBK8DnHODT2pYeDlJgwM5YQ/NayLGFLosWr0aO+VmhmvKUFKWHdmy49NseypMSoWDTq/nD
2iqxseVt8+svL6B1RiQp4vhxn+Xa0t9OYeXBnaII5HiEhmRNb4w51RLZNhri/BwdgSGf0LhPVUA8
i1QF16Ru8V4JB9nXxGivGbsv5NwN9H45m+LnR73tPcKaaVP4CT3ez0zOB2Uaj2UoGoNaLYKtV9eh
zWTMhfEU42LQWEk68iFwV4m1P6jWUt53NZwS1Nkbz09qZvs/T5GvSNVMKob9VnpR4x0ZhzsQLGaj
2zKgfcRo/aunLEbYeazfDBt1orOl+4YilzTXIK3Ea+8FPU4OnVazNNybzj8E5oK558rnwDAdlVl/
rXIcp0W9uxCh28zHPMDVLsfnnf7jD2yyh0gC/GtIHue+AaFmtoy9inz6ju1HUGGci06uXfptpyqb
M5p1yeCqDzhISTNZR6qvSi9ktmAtM1eOzFzdLpwgbZDbmLsnJlOcbvGt4UFUKg3iO6XsHns5MnZG
+ShE5/h9gTD2Zm6xRe9Uqq2E5jzqNxIca2Tx5UbJokTKOiC29DxxyrQ7KMBWshb9NWTdxhgHOH/O
1FKkxbdFqAdD0M9GI1S143iGABtfuYMSKvUS/dSQkdu0MB6oTOl6Edcj5yW7YILrSNs1Llw/eZrL
0tBlsHK9lS2/xHmvtPqPcMptNRjfjj6DLXbrQxcJb2OedmE7ii/hkJYFbOFZZ8DisAjVOXWfXfEw
mkGXhP6V+HV+pIz3VKBfNZ08R3m4kBugifCJw7yfARg8Fn0/uv3xxyFK9ZvNg1SE2DRpAMc4WF2B
QKIj9aXeesYtVT3V7TSXveavn0+Ja8GlW6tH1tf1rKLwCEboi3QPMS4z/Lefd075zgStzkKzy7Tg
rd8NEXZ8xhGZa1uGKVGqnEHUUMp5+bDT/RBpGD0N8YCYpfrQlDBUYBKr3EQve9D8YUe/Z9PiiiS0
n7ZYOH7vqpU0LlmQbWEAAZA15dhd3sD+TISQL6mqTa5WOAHLEL9V3P9aigPLmRHw0LmIvU+0L11W
4SlX6zwOTLaSDRX8z2kVR10xWCmhJIRyiECxKqWwwOv5U3wxcsavU0PvM7ej4rOzZq+jBLZB4cm/
swZ044gHEvxUUoDt07byC/KZ/kePAwGzchLOjgR0Af0epblqiY0kSXkA2XLc34r1fuIZ5I40H4DM
qjkIumSqeWk3KdGZncuux3151lu+JQ++HXQ6ysjRHyvfLKASXqO0m7r93S71kyzBKODA39yJ2RaB
NQ191KqM+IzTtOLRnHtffKkHtSUzu1kWeU8ugYSP1TqrDJuFJWp5NtUbbulZ52fyI0TnHjs8g7T/
DdxTmfOl4KOxhC23oc9yK++E7Kb4DeBBvh5T/SSuIpJS7+mb1A51hmqqIBNbegTHFe+1mMAYHfqE
3giJhBoxzo2RXAQ0ejbqP66BC1q+SGwgbn0hye6bUxJKmKc9eWxbG7Y2gOvrWZt50SqJHotznX3+
I9iAGi1XX2S8stNITuuhfX6izX33InU5O/TlFwbgEEv12bMDt2DNHPC2ywQWhZfo08O7jODwLW9B
Yox28z8EFHOxcOyNlALjdzoR3XY/joZbtE+NiwSPEnA7Y8I2xtrcXfEIsmWffxUpZqEJ9T86BRvk
wa/lSpHznr81FAqopL6qZGWW79e4m6g2VQBTnDNFz/aHC22fWfWpNZvL0/6u79H5Z3m3a8xFhe6s
hpEdv2p7FTC/7OxYjsEHD2/YAyTDLvugBiGLSnMYY++Huur5htU++L+GGJBiQHs1Aukajr32p1R+
MJXLwpwF9S9kxYXWxAE3/XjQQIbli5o0CWNPPi0w3k39zml1hfRZzRjS8ztBjpZs7wCJfaqJF8tz
k/0KpYjU+p+IbFvfL/yG/OIu1Sqz21a8+9MWtcU/x2q/spF7NlLxruQKMtsH/hUiHaIK5UDhHJWZ
9MRhiJvMFMF/tij5lb2QK++uJLUBEc2Q0MiPVI53tAfUj2Rs11NhfaFrxNx+HsCp6RftkkcKCD+I
1L+5TA5aa8LeSU/5VqJn9WhTPoU8pdPK08gzPtV92D9GsAHe0XYiXDZm+8tv76QH8RZAYQt2EtFD
+BFPalX9TIa6q7baDk/FdtyNgx3sSBn/7+y2DlPtXr9qnn0pAA/+ZwGYosNUxy8xkhI/V14GE9QE
xxtaMtbF+fDlUOCAOMQwDXZWvDgDe3AvADmo8TQ0x3bfsU7/IX1u9/gkgqPLYvD4b8r5DYyqXpOr
JLMNhgvuyoxg86LQVC/DUV6fxhP8kv9eahmoTqZ3+PeWy4Zd8IopVleaIu+zaEAMXx7/iGd9wDMe
xe03lVQJdnSnNein4UpFz7qxRplJ+rrfHRSjS1ckrb9tSawGGIxId9gL9gam5rEWld6c6Z7MF6Q4
fDLp5UWYUzASuf58zNpJwOo6yiLAgAn2b2wTvaop78mKvnt5m6KJwwLIjpM9TxVAuN0zbJprjzJK
o+qCdJQ9ImzsEbud8zaykTg4/d7nL1TCrLB6OUUeyPFYUSsRHDM7PG2pI49uv2iZqAZJtG7zKrW6
6MwtznkN4dvUtukSswrXoRkfDVuFloy0auj+U0eLF1WKhUumDtItqaZGv0RVpgBUfMpX3SCBbnDc
O5OcMrqttQRU3w9sr5bWgPICSZ1+oleV7X9SBqHRAtytfofPMbfblJMfeBPwZRH9Ie5II7ip1NGr
6ToomMu4FejKObwwvhe2TkTprCmfDavf0NOyBncAkDGUc9fmkCWcVCohrTfmkIdlWf2jKHdIj6UG
RYz5bWyUwnmEBB/ez8xQJ52qIOxucqHFR7+O9Ann4ITYLw95/oeBYYrQV2+ATCx9D1UHrSWOGjO9
7Yp0WYu/jV4kbzDTTonFph7Yc1z3EjdsmmOsDjDdvXljL4HHZSMcQhQTWPLpf5SOvNJ5ACvpm2Ed
a+pCurYmtG8zF9ysl5zOJ4sOOX//9uyCxlW/t0rlkkT5Z1qRfn+yPjNJhEfw0C2WC5TvcXbshTbd
s7l8xTpaMbKAAHNYu6R4o2UHfnlvrFFsU1srsOm2ut6aTbCZju6Vx5PPrwB6/Bil5fkFDo/sir3p
ip+oQMvlSz9FcShMZ8e+l+pIM0G7tqwpXxvtmgPEQtneCAHqLJBHinpLQr5jWhlp/6AGwOM+bb1t
lodoQoaqw7L0OchA4jcIyuDGZSDfD+HRoSUhN9lezgB5nftZ1FGA6puwxFeqkgziDKiDIF0bVEF+
iqqFgtwv7aKNaL/BiiNOp3w9uzlx/+W0JyvNKV9C0mN/Re0AFUz05TloEC6KeS9fK0p3NkweQUY+
s5grsTZHxU2asba5cW2ljjeJIwOT260DP0Hw25jwIunsZD8c3xwrYQ5c8O0TDaDhrGfOOtgrJKSJ
LWGpKUMWX3lUVHN0ElSOjuyqe03GemxSAvaPlP3GAJVk/md4sBXcUhI6YABw/kjVVzqYKy9dWmgh
ieJvDmpX47gslNcx1DkDBnz8G7VcEXmJu9mSUaD92e15/AmcQBnYcaEZ8Nyl1K8xrSctlykwRXbN
XNbdL/8R8LH0Os7kjaoaxQkVjbmczHhvY5moO9nD7a1yGz7mecoI2ohQj64AurSK0PyjwzqRg1Kw
kpV/1muBbXoWy8DaMsWJ2MFGnzlZRajwXx49dKBsWybBkTsnqqXucxzrFv8jWYaFijHtdw70/6LZ
AYH26cDj4s8WSPgb8/TOY5x73ls2aFtBBf5FQd7i0BDios2sCtfvwnwy0YEc2ImBQTQDZJMd4OsI
k9z90+F2aUxVw1b7q77b8Dkg8LFkJyRKnIlBhU0tfmNETCRdZBQsCNJ7RkOCuIwPUh7ULu+XB2Ll
xaQv/+l6LXSedpNexYMaYUGnNuOovsHdSxgBXpD6ke5V5eOas9luyh55cq/u8Q3j5zJ4H+PLNfmC
6WTsa+LjFVqjphgSAJqmOdJHWcWiFoS6HbURU8ygLoeORW5viC2GRkbQ9JL8TKdxGloCPINhkz4h
qqRljisTkBgMoJIo2wlLMA1FNXHbx3eyAmnGe9FHRVYfKWHBdVB1FnMaqn5dWowy/QPrH4AAfwS+
aYVyhciY/u9K4Fru8LRLwS0tGqfgfvPpLNuXOZOT+bJY+RYCiqibkGPTzS5j8C/dusfDWGlvNN9l
E5UW6DN1V4KXZOJI3LRh4+cpjyza98sga/A96cRJh8lCttpzKk4EQMbUSYIPtaDq/x6ehlFvEMn8
FHvuof0YnNz/VxNzYqguxwHm/vE2ZwQif5DroKKtt4Eehr5ItYA6VNDD48fC/R+pbRRHiiyoybHC
NNQJDd2ZEGADoXN/DpzUwETqm9YXJh+jX1nstwffzn6CF3cUnE4GSs6dOUvFM5ryEtxw3eQb9Flb
3aL96CnHF1x4v0sHxLNwKFRN7IlqwLm3w0fsTfM1wlZdn03ssuEMKffHIwIzY7wG7pz8dRGyk+5K
d7Ox90rgschYBucrzVhdYUhfW7yaaSGe5j7sBNJ1m6/vr6X04ggCWgqi0WlL9sF9+LBk4Jud7J8c
1LN6SqJ04fHoWQMBBK/cR/TJmAyPBDA66xlP+7JYYp8YTJ0sAkYiczaH5jBupeJ6yiM0Z/0v+VTS
gqjd/sBXsesd32PDxC/mGphCJbfZ4Gyp+Uov3xN7Y7xz1fGwH/b80ZCDW7kFsg2uyY2xHpy6opuQ
kVtxonkXWNbk+lWE92/AZDcEhE6mWtvRF+J4Qj4E8bB7o39z7NUlNF+mfEhnagc9DX/NFTWeNkMf
+Hueg9DI/UqgHjQ6Ig9U8hQVK9g/+AK++ffA58+uev0unYRXGRvE1bd4fMe3dbAlWCsRn7NflPkV
wHBMnWQTLuh2lJHHSiale567oljW0kbtqpQozI0gFpvSAMXEW1ZoZcvk0XkkmYTaq/QnTFskUWIV
n9j3bVT/KTehOgPos+iMff7FLwzavDqrM1mljUU7TsGK/Qon41aG0DVF2WegtLH8JTvqd91JH1iC
Rr1CSqmUbEJd7oW+1u6RVOedBLrX5bkegUC8Xade2MW8E/dTsrF4dkqFvfAzyrzj9gW5LtV5rx69
+5a7yNQIdDs8+HAcQ7aIv4D1axwQZX+oMIDUmm9Scf2wKkiP4VLuLer8zkoDTC23lgzIP26rpYi8
xRUaVz7lSkR7uyJfAprIwlZCWGBhGe/KBmYhuB4tso5M/R91XIamFwFDtVf3KLlceavOEv7vu83s
jfl/aecZNjR9jmVE+wdCOmjYZIc/ITE1ss9RNiRjGOsbEItJH0jYtpprYSZKnFS0rsAyH/joMtQc
Wd73VgC/yKn9SinoiOCJG3f6hItlYLJPYh6Oci3l3yTKLrimbRaqSWgNfrzEQC60Uuc2y9HDe9z+
p2Z6gWRxA9MNMJ1UvAwBM7Lrpr3zRiKpIdxXO6wkvPxhHMZZEKy9FDRv7MbjeAJ6ao+fNuxRsXup
dTX8DAosbczir/vfdpbCjpo1bBe89Kv9AsFcpSoEP3a7gyZo99yVSK8WpHdIKY9KRJXY9a12Z59a
bOQ8fOuQp2fpuWuL9Z7r7/WoXcvDX3SlrQormIxKbuv0sdALd+LIlw5R5zl7ZomwNCvicUdSXAqW
lgEP6IeuYrKpjrQuWBhei27gwygA8vIC5aIxP0EZnOltkpEnxDIlEzLJxjRibplMqXESTZ0/UwG0
dIonD+gUpI6Z3t2OFmLKbfxNF8ITEYguNFRqBBkO1afHuTIh02EtlLVhAMiz711jxJyEmXg2qahf
BWQH8zllgg2xFp00+YaRg3IHCiUtnQCgFbIGGwd6HMAjDnVx06Foy7CaoZQVRcdmYfK7ONorSinT
VHPSO7ngUW+12a4fB925dXu5i17bQt5u6nW7+gwvCcTkHTqXl177FfS6xZUSaHjCFShSIuoQEIV1
dCqQ6HhyCC2/lONHqvzuDnFUOLJACqCU0YI14oT7VglUaZsk1dPpjM/XhAGEl+ISc/jQUNRXWAZm
UnkCPl/Zi59JOAJvpZHW5x5oToMZF1Vd+mVioNSZ8oPnb2REJ64Fs07XQww2KcKrYAf+LhNcK+yz
6W64QmK6XmjK/Jm26O4mVvXYxnrjc5aMx4yItx4Vto89pOBvXDdCCPCmLQQlu30OExksJ4pLRkes
UvEUtXrcGU4cbR0MXjvQDizI8xy5lKKKIAEiRgwI8jV5qSH+cqAqv5I/+1zUaDCOD0z2CDJh4ti0
g5ez3DXxPm6F/aSyl6teycBdGQoZgf8LP3uIgqrz/GewriwCBmGl12WCYUBiUzCpVPfnvq5wgCF8
rycDJZUl4zXjfKRHozlicSvFn6HUkD2v/eCUM8rYbr6wOT0IxIsRuRqbYLohVcOwWWYIJqgPElLT
FqTwCiz9/2TfTVupmlK6CdpLNjYa4tb+m2sNUZQ0ApO4wHNDuwi2QRCRrntf/2wMK9EsbmbrYknF
QkMk7t6mv/MbODUrCzewfdFBmmwtLKCPxbRfe7C7nUedDlHR45DmTHh+m5CtOzkxIoxOYuUReUp7
7zs6aCZaNMR221LHMuQZBQiseHCKL0o4uozed1mxoBTgiiPkMgvcUkQ9BoRPfO4F00D/zkdRcOz6
7YzALbJAumYCREp4pc+kJJxLRgb0sxXam9hUo904GaA7DbtHvbzy4ajIL+ZD3BGLv1WLP0DUUvux
AqKZFSlh2ZJ6UUrasl7HOqWEg1OIoHrhVZ1UBuRtyag/Fno8fUto7ZPvSMQ9XoLfxc0K5vQ4+/9a
6ANMsEP79kHOJCF6LjgaGyGyBSRzPBjy7BRoNh/POGIKVPhXmoTBb/NdcWJ/QmWB/3soLDvrVxIc
xS2aktZeZv/bNktL2TqLiyqrRVw7uwLy6FibkKmvlKlVoiP/l6C5vgzMbvz9WHrZaJ55jym/CIT4
iVfCNFDOWaa6/iMguDKVzGkjMbYNxSdyTrprkS11BLCuP5FKrwSReqBBNq2eicSEDWgzTzhUJRGT
I6VvciH9M6GKaGHEA8KVlAxGZdDQpUfFoMmrbJar7dAd7p3LE4G6HgWasn7lSK+P75ZF6mRLi+Kw
zPlSBFXYMWEXP+/YhGEiMFG222cx/RFtOWdsee8/Pr5NWC0KlHgZA++x1AhgT5v2HAeuJvhKlOy5
U7l7slVtK/2e/G5Rjh2dXWqmribtM4/sHzEOITb395gAVH5mEho895VLKpWec7rCPJEF+I5yZAcj
B1Xc6djleS+bu8de2d1Cx9etSHsUA4FtIBDpFbKb4SXIqWk735fqCAUqyXFTajgtmFcP1i49+OwA
QqNuEPtk4khLxViNgs2g2dsNyb0TdjFTD3RcljXrEqVi/oNJQqylbcEYB4b6nnaB4lKuGuhJ9uZt
PCZF1hrzTc4Xalc2O30LJ8W4fSVchmOAndWQGOAokPWsESGCoeBq+KbYlL/BN+5wDDdeA9v3dPF6
86ZIcxzm4Xxbgma7Yn0DpRaF588S0mdnrOE8/HqyZY5Jvd1A+H/kCFnwcWVCgWoQBW55/ObxYMFy
/uH126A8OvakVfZMhPh7tRAKdJsedWyAQk/igxs43s3j91aAA3tSyp+8/QtanQwDF5R4/MdOnVgO
x6vkKvpjNXbPbM5dhwfN+sobSOuOOE4NpMcOLZqOMW6eoDbEFRT0pqmA7H4ACC/4lbTIuB9E8BEJ
Ec06A24+VyO3rkAhuf8mX6jzNkBx489xnXflTxQFPtYZosyrigFJ96UiKw6Z7eGUdCGwCc6juBqY
HfhZ1J1i70/DF+WabezFsNTO1p2cXVn8PiVJEsdrQR6QQEmzt8fUcdtM3FJs643WvRhObTXWLSba
mukSZ/8dW5FjQZVx5rgYCdzs7RD9bL2aTw1AhaTUsggfF1g34pvR33+VFfiEawLcQ0/NrG+ykPkh
bF2CGzXXjeqMfVhw0YkfRHzUuJzEvIkeTx/GQejApWiLLkPsKHQS31IyNoSSwt0PVxcX7QTKd+fH
BmD5aJMoPsjjVWSuiqoU/Aqgrhj4mBOwlRcyDkqQyLPZGj3wG17JWAicA0NiEfXxTravUVzrfy/f
Ya1GE+RZ9SO7S7moDl+Z5lrY7o3tr/csO+cLQhixZRkqYybaBpO0sU3mF+XabvixKefxq/8uWQIO
dxwLLXQ5yF+Dogq23k76x+YtuHjDdShLSKHFr4Dv3Q16v3JX0ZFCgz2fH/bJxIZEV7EXBaIPxVoy
pk3ylRqVQes7k5k4CkHiL98SAQNCgbbxYJnVh+NcyKrGUvDKUOZ5g8vJ98qnABRWfLElXcS644Hj
5Qm+a4QMlL09gJUQMogSQKEUFzMdGTNLjw4V0rWQrQxUxnMBX1nnSsp7QcflO5tKkT3rJU56ivDn
olO8hMU5ChAF38zVK3EvDPocPOPKA0aYOiroXdREn41zT/wpRnjJv/tZI9zIQswUsceYVwzYRPCT
Oy+xxy2OIQ/PvF3LvpjUAeC+wSepAyPM00vJ631Yen1mvt3f2jYt8hUfAe0l8y+Kr4odYF2sxPOO
TtrpTnQITI9Zd2MpjINX4D0OV02bvljlshPzyJ2ApAaxl0QVbi2RysusD2jCBsl8Ptzg8wt3h3Es
47CbEnpYrF9OBTOKXHtitPGLi766bDHFnptSMZLSoBN0zf4A7ptq9CvrtNc4IXUitCxUZ88W1zEh
Gz4m6SnsdNZtXRPdEt8MHN9GeG98DrVZ8+L386cS6Av4F0axCV089w3Wz6fe+3nuSEh/bSGjCUKG
Sh6V3WXYBC+w2ObEakr0s0pfOj8crC6/eu5Yo3dcqNTUBocf2X5qysVjt5wfaK31Frw2XP/ldrpf
OIHu6wzTn8YTYRhzt5yjSwfVPRtac/s74x+GOgivWtEgDWXsc6rdL7fz8GnH1AaiUHiql6Jst1vw
R5ZdPDwJrVnMKNgWS5CaX7ru+tPVQ9eY+yOO4/vhVGZCfs9+cQj6qq8FzxAELWrLXN58GPITeBzO
VPwxLu2FcOZ674oWlrHs6EkSR6waJUN4N/6EgSmtMgU3QCFw8kiNXq3EfEijVfb+lKJ9xWUXu09i
PFAuewong5pexslGfQ8C1B4lFIP4dfgFqKHUw2kYoUOe07wc+khBrFZzNNsQ1Bs2kgOrMaA31ucK
vmmuIvFz6NGxgbh6g3ZK0Qp0qxu+ivJO3zvQiyIREqLCg12lp6EOtAMbbhBUl6ZlplVZi0jOefRT
+X39i5jIw1UHyIR67u9p3Vj7cZKwWrS9eLXvw/3HLDBFwNvuqXBF0zicFMvGtwDAoF2gqXjAPySH
tQRQVn0qkqUiqfawWXLkAd2GGu5OnIx0Ce+KPVC3Pt8cl6+1hJb2mNBjDvw56DlNn97q4p8wNTLz
JNKFEMwYx3silgeoByDS4mbf8JMHoLDyT+ti1JCUu5SEL9SpDJWkzMOP3pO3EFAMt5fjjtR1l/tv
wre3E+NPndlJOVQFW5KPUTXuUbAYFVeeFUERh0eKsc5kUFN0r/Uj5UMOmreT+TAohos07f/FZzQJ
bQsgMeABchgB5iL7FgrJ4pF8BU485HwclXOJYsi6hUcThR2csY/g8IutDFrojnoX2lw1vx3H/uEn
/pN749ypwjGvg3i9vajEdeHFS6o//u2FH8yJONlCZ5rxcXNIBtzp+euyrSoXhum44t0QjEDB0KZT
BPwdyZWWpANguofqnQM+Kic8vsS5Y9JZNzxb4COp9WcWRqqSzQrG0ixUVbszz3y+mef+2l3cFoXz
wXvz62y4aAla0FNMe1uWgsAiTGx3vqg4RaBQKTwZf/dy8xjOdTL6s1Bv3o1bT/absQD7eD9DjP+C
OvD0qwDXn7u2W0kCXqs7XOjxkj7+pVBhB7WuGh/5RYacJV1G8WbSuDhxsQTyTaSQIRvja4FuFleD
PAE2x4BnPKGyDC9ftw3C9bpyTAq7uXViulEUqkAW7JaM3nat7GsvHr+/V52gMqoUuH9+Q5uoX07y
mdrjsAQ9RawEJ8LuNUCCWUKWjuDjVcj2uEcwG/yglKhbrzJx6S66jqqAly7nYB9xuxJXjWVInY70
DoagZNERts7ZqissQ8qBAqsr1ta5gwCNWLuNPmEbSzPNKpzgEmKJhPuLSfOJMZ1xP7zF55oVr5iu
C4Tw73sMOZaXgfZAftA36836TtcKan4D28VR8MLG/hpPeqfYSCv6vHeiTS3aFxKKCgTf4tRC+510
sBDwoAVN92/pjKanDvIsyINuZt0WYUwxCgBLTEgDI2AImcrlCVm5F3MBTA82mBeEWSeXH8yGj7zJ
NBaXcdbfmW0Ktzcw/ZfPGCg8Dnay0iHfIP2qwcZi+skznJnFVFgiT+fQaUMc/ZIqF64XQ33Em+m0
UA8TnLXQ4X019NPNKOWe12EwasL4hl1ZTP4prvplR9DVl+KA28ynBKhk55P20CwFJprgu6lfnjIQ
nNOmhDcoT+L1VB9bQddSWn2IXPNSmM3CXJv7bwkKJnGElWfMdL282UfC6iPcAEw/vnlvN9uuQSgm
T2oO+2fjf8zBRJa7rYLcjaUxgKuKIQwWM/0QR2VGSXFkdU17mJUgjBPHo7sM5EtUrtcdQQVFC2qG
cy8swfB6Zi00pOpT67wfvVvDVM6HjrUcJgaVSgyl50AbWJin0onlOXTLfK4gxDPtabhgb58Wu9Z6
6crm14rKwpjXlF8Ddsmy/bhI+MDmELxf6OmvdBZKrYdFyWEDHGXYB/BOuqGcnR/dyZID05t3ixuo
IfxwWQjhvSC8SL1GOfDQ+Jjdt0ovqlFv0qM3Tp5W/ol4eZUcFsKM2yWWX09xzeY1gTlpaYMFhues
lCKKz1BTe+WuAXjMfX1vPXN310Jnnmyzspo5sd5GBrsYSGTBVwQ/CYpNkSFVPGHLMslKSNFpQUmK
jpLwJdFn5A1NVLv5CmXeqOVBvJkYzTV7j4lSeL5SE+cDuWTHaC7c88vxKHshERQ8UqkPyq+3Zbgh
RomSOxCuOSq/LqqPl8sB5tyHLNxhwCmmjObWtv54/srurbhpU1D0UJ+nWqwNKhfhYlr6zYgx1A2Z
C5uDF+dTb7q/cc6CUC0kIub1m9Uwr7Q8CfdV6r3jg5WFsyFK1xIzC1yfoXfdbcnt/7EiChWVQ7Jt
iplvwaLZqAinTJGDjzlY0o0xJPpTGbicD8kPZYRbXbLzXzMkFE/bhaeR3TJeBOv/3kk3woIF+xxB
Or91+j5/Nlb/D5gi6QliLDyKLXgZiucED4SmBCcBswXSjo9r7joA31eSa57h4d7SEuL1QLXJdCE8
VPdVZthUVL6d7ySwCuxfZAs1i3A/9KX7MbfpwxaCDHbCi7LNdOFuQCbyfqn1170TNG3cvXoBbBah
HsZkOKzofwk9p9EChj5S7/rZFQRO81r3WCvic6KLJi4+WY6Mh0dDUehc//1dhjutqAPQyOEPsvAI
NeqzcAbPNC3XQwQyVmmmmvy4yRw6YUeIZlLc8B9xx7zX96TM0AcHWMAqosmuGzaXgvnuTxW/7Yw9
f/rqhJEemGM6QLNvdA6715dzvQqqdx3NTew1tk+bCTs5TsWvWPIgnKadzt4E69voq6q5XMPKfQmc
5u8ktuB+DgAMCYAsRLRTv/HEVTidRLU20aXZtLtuzwZO1VWeiYty9pnItG6H3CXORyB6pfXWOFwP
IAJkOzsq8mKcdicgGhzPdTbg2k+HSCcraj3es3rzD8hksw/tWdY4U1VbYlNTmHvkD/mhyO3NvKb8
84gq7Tx37m/EgSkkz0s5W26ViVjeeU45WatiUFvhT3ZhD3HxUq9XQ5nFiHVBGMHNgTUNrV6MqeyG
X38OvVmWx82oMJCACcAdRm95FxbBfEPydbXBG/ZZiTIILSoeABVoDvqgpvpHLF6lY0GWp0FZMHI8
IfMVZ5Y3/FTmaq4QAOxQa4X2GP/NeSPDcDCgrqupvbvHuAC81wC9aAxURDMf1TXs64tvioYvz3AW
6sCEkXxnRVeNdZvxplXvKnCyXkWlfOxTB3NdBsB5Is8zDJK93TUfXq/zAz8ZBUnhfbnJ/a7L7CaY
F7tly3I2A7skZMkVOm556A6ozMjdEa/slwQr8M6woAnn9KDwl0PqMrn4lUSN+bvjzMdlx6+ENVyH
YUOnQPVu5hyWtQxmqZYIf7Ln3IYW3y1dqkFyyUqPu3XlKFxnsc9Ft7fiuh3xXEr0HmGwfgaPG63C
0f6d/bjs85qMcbu7P/UzKeFdVADIZsxtwX97IClodI5YAaVItYTlNh3KdqPiq3msa9zs1B4zXpCt
tIXfX0SMMDXX6RujFlUHej08WMS3ofLp5kW9qjNXuq46AAp+KzxRh/ZPVo5A4id5G2GI1vHr30/v
tzSCiCB4VrUqtgL1lcsoFeqDmJ0NYB/E6RhZeBJmeySa57aV/TEidpFTgglpATsjMdKAVfjBUCAM
FUo+vw5tkIEMxM9TjS6hnul//whkcrwpKfB59xT0UnfX/J3x9VFZksoZIMUqYAW301t5M70zJVtp
XtY1RyiB4a3jXTflfkBS7PXapIPLVuzJqLUTjDaLWxaXe37yOuYmL/Z5mvm0/CY2YSHVhAIyML+M
5HIK3MI2L7WvoqS8wKgSqWgqEnYI7xnwqkMcGyisrgu6eoGYOgdvYpnWBSZBxz6ecoQe52cLxtsO
kyCQKdkv+qwpJ4TqoKEH+lm+ZO9K0XxUd8ZPDwUtlz79pMlgIx+OYG+SotbmTzlE+PgkZULaMLuy
Xo1DGkOXDDowa1CSs5oNo+R3pPpfA9Mo0kDAngt/4gyls64RHS9pQWxm/eRb2F7ycse6+YxRE4Nh
vPdSxHoLkrROnWTE02zHd5yKiuQ02q8MW0U0JMoedWZYrlkAEwp/cgFhhC73DhENY+fiCXQ0eZaH
ZCbEzLnG4InelS7zqlF0Tway+MZh/RkSLqW6uB7L98/I2thAuUIT5NIDg4ntvZ5cLkfC0IXRs46Y
hEhzB8ilYoIQYKZxMcAGWJ8wP9keVOkOnENK9Tu2TMaPEzI4DSZULH3cHtVP5ykQ+lCzpfrK7nc9
6xdcYCoP1ZAs8FiAd8m92dslFYZTUzMCzbyFUglu/pxFoOuJugZYtblQ5sW9J8w82NkiVkuBugKd
g8g8xzUpgGMN6fuQdcl/yaN/beoZ3rtaNlL1pE3N4OxhiyfP6eFuxe/XpFo47XrN8Pgs8b2ELzu/
mL9oxzW8eQuCSpViDNG1a3ctoOxLztiXDEHRc0InzVtjsZz9zrmny1aS7zh1OKzJQdWDjGPLKucT
OBNy/c2TgHauYYJFQkWBOe3yGybYRUH8y2TVuIvkUkL64usDDDhFemLXhMSnXJgk/at04IjGBBSo
41udY8Xjn97Gm9H7fOlJXLzBuDR6GfYSjFqV2vDN+Gp8YmOMZO10s117Mu6djlH2Tia020aUHhzi
EbJhGLz9Tx33whbWRw6BxYRj/BOQm1HH4kCnSSCb01HWc9FAWVuK1s/BjtPPZ7jEMubyZhfqFCPQ
ueX9ga++EM/YBacFTGCjUUrQm4EuqsD8KKnFZxlUa+id2KfCkBrAyIvHUHTRKOGNKRUW3sF70KdM
NqqCUOwU0E8faA54Q6HWR1/9dE4tegYn44F/2kYilYRQjScI8FA51OsmXktxmVSfkiiIcHfWnGum
CEOBJlOhxvRKn7D/tMsqyhRWLZuUJusIfH95ExAEg6qkyG+l3eSllmapYoR8vGw39n7V2v1WZYZ2
5h87KRFtT6f6Yrd+BveIFkfU4l3ZsjUOyy3SGJobKBR48/KJafw9mbEXOL9en1uLbJvGDEOJ3qN5
zLwU4X26mc8MeyYgOkx9k7LJJa2zk+pibr96H4sRHqVrlCTYX0AIczPZnoqoHvXRLN/aLzoANPNS
V1K1G0va4S632YYHYjKhmJh+LRQdO9GneWVJ6vt9M7/S6ZvFu+GEm/PwgYTDHI8yrVaeUqjiSDYi
hR3YGx0uqnGEA85MxUD8/RqFiErHImKbdmkM0y/eVmkU+qCNSxbLk/pEZ+F/IZz/NfmnD7ILcCYL
6OK5iTqSnXHYqNPG6BxRqVEvvGgyoFPfMHkT3Kw0mok56+f+kaOj/QMOnhKhEcJb7Hq4VtINfsl4
91cCRAjdnbC6DLD8sBbaLbYjzxsI/bFb+by00xZUlfKuxc7pnCzqjkuAaqtex8J/h9QHENPwO+Bw
rFjlOgK6/bD3OcJxti1v82NBKmlRF1XvW6HKuAJnyqdaVl8f83dlwnXgUyFfb1DLHnrzUUkEMPCI
4dYFVua7/ZvzD9XmffbaRhFh56/AZ/n6I1M5Lx7t73ecqjzxTve6z+cp1xSg1hxm5BmtqUe0LB9t
f0cVcb5S/6Mh5n4j1Fpc1efE0iJOgiVYqCGUk+1dsYGphr/zPlme4hIQ7xV/7iVAe9Aw4ZzafLQ+
BnCWax2fJr41tdVpFOcv5WSqta9ipn8bl44e6HybFYKHlT9WhNJRCH1HTxkkM//XxYSMe6jjpTj1
p763WYAkptA+YPOak+VgSBofebl8cZ9bhxPILUqqFyWHbovitjIA2WaaeIrj5wWJQ391BH08VJ3b
CX4QUpEKtis7YpiH5jhx8EWCS+3M1BsW8seW/sJyiijslvZ5O28vA9WUdJetstd52TLR6BDBD0xx
qkuargLLtBJDJcQjv+mIaDe94smSvsNf01Yfq2qi9zBwVFgQ6gyU05mjbO3h5myJKojlqAgaf0rY
SubdvKcs9LW9wY/kYhT6g7f5gO3ysxl82zMToyM7DaTLi1FC/NGNpFAg8STQcU1gblc5dPaQBikf
40OmIo4vCYZSm1wrrLUGat6XCiK8AOijZeF1qy9BwFozc1427x9yOR2X8fooOcd3/alS5ubJruGT
52//cDaPRMwqGrrWQWv3+saz0Ohc1Pbf2FK7Yu0pOm2bslbJ1516ZxEJ9K5F3PuDKZe/Epkjl2VI
FfBW7pVRBk5lMEsBsIbEY2FBF02UQm2oUbSHirqqwIrceyY2mCHTuhxghvEMXaRtOidfvba7Cp2t
9mt6zqDUyTzeVqa9vzdQLgf9B9d+cnkUFA53rRg/rraElG8P+WGdLVYLwfk1F+GMRWEhtcdAiK/N
86H6SUlJKPWOfQgMtqWTz7zQf7mjnC8SFZFPk4KV7wI5Ai7JZQ7NWqBOcLqSZK4wJlEgLs7BpL6E
izqfwueeOkL1QYFrBVJJH6qTIT8K025qrQySBGoG9wbVTPQrkrCfm24MwIQp3utZowkl8ReBNTTy
rnbbhhjI76z0Dm5fxkCYHWR8tt1GVEenVI6AIfUmFeAnovEPmToql1mXmmjh/IafH4pX/LCvujJp
OfsYiQOro2gMm1TK3mq+F9ntFP6bfd4sXTLjaNaCkJ/y9gmEpC40cnjNxeVfxuYumoGbIY7omzvG
tNyPMVF0kzzG8lKxKu+BI4WJQ2gqPC5v2m33aS9dv0V1disdUSEsGMYqPjQwTLwe5RTvyeQP9HsX
vOg1cqH29GU/oOB8tDYI+OkIG+LgozHUj/5zLzFx3SacKNCxJ0dEo+kfbx3C9GjV8AEhQuexrWgO
pZJiL1xfqRROY7jzYRJ3oKdUsy+ZWt1m71H7vRDbnS8VohKCcDS5AYYUFLcUjJNK8x2SH2nxoEo2
AZ6gZvEjpi1N3Vg8WoXjty96ciy0fm/NwMRhrVG5YtTntrVEd5Cmpz1mN2woKsxUjIozl32Vcpgm
7uDnH3nY3AGONtlf40yLnDus88SMerCyqoxFfZSPn65+A0tfQJ7vLl3ebyw/CHdJxRPkEqqrcxnc
m0+nShRzylF4hES6vfrWaPEHQoT0knyYETJNt7FjO1FbCWVmn6Z2D8AEVqHUs+yx4MIFAjJy16cz
E0sHxIWu/c6xzgXqi8G6kHDKpkHLexaGF5ogN+tUzJq4TKNMznzWK7Hpn221lW/dt/p9UH+dKMpj
jtVKzEXpM7RbOk+VD+YM+lXD9m9DN/eTdt25AJtXlOKw6yMqKYYVDCHmb3KLtkKQ8j8yK96Jo+ZC
8az4GzR6/zQ5WjD0LFu/fsWBIpNy8Rr534KY8t9FKgArGa4hXLCAkYumH08/0jCn5RYX1iAa7fJQ
BpZDDfC1lOFCDIRiRWgyasK9E65oH/p+t5lVI3KQFDRUZ0F345NUad0vmTVteG5jGkyUry27LWnl
Lr7jAe9R3/ZH3pTmiLp6csm36cL78gUfsu+tvcmgozD1EqUtmhcYPsbAUx+0jRmxia0mdMwqHShL
uMaeSa1b13hyiK8LY5xsuhATpUDJ52X7DE4wckTgvEgnrm8m8mCWvL/WBkBnkLZzHADTaNigcLfe
UMvEn55a916Tn9/EPJrwL3lRAemlxZYzQhe5NXNXCjBGmsk1lgEYx4Pj5jKltS2FOs0oLgoYeR78
IzxDz7AbFQddZZv9rVxUUMNqsP4jxSXhgFJZjHlOPG+Yx5GxGSomjF2OwmslSrG7wamMSamvEb4w
30T6N43I5axZhg8uhHcVUbqis5EaGjuIaAbKLn2pV/cAqXjbus7u1OBS2Bs6EZNasDLzOFhEy7Nc
HMm7IalCUCAMtAtSD6rQ+UJnopejmKhLECH4cA5olUaX/dZf6sEjCDfBKiDZ7lqYeALkEKnl1yvM
SvPbU9reVjii4IwmyFYPvAIJ9+oSUpB3fIcmS52OBDtyP4rnHvBpjzEWKuSszbacJnklpkIpEqiV
exazd5sCxefoKPnsUSQtfl0U8xvXiASaL0mbSjKhMIIBZyUyJmxYyZAxs87tz6Jfp48mktKn+4Mc
TCOHbXP+6qbOugARYQxfrXN14Lm/1N1//42YRAhhqxZVmFInMnKmLx9tTFvbEVn9p/e7AR2sWKuJ
+2kTr00Xlb0bV1sssJVd7QrZ82p1E5dfQs8LqihFMU3xH8ldFDPu2c1znVzw9b9EVL8YPNw94m39
ey2zVc6jpfXSsYNrCJebY6/EOFxlhvhcwb/OCbQc6iRhSjXHXpeOS8XdYdm1xu1pCYiPtqr9yepR
CszTgsABX6dkFMUDm2tSEL39ETvTz9oFhP1HWxbqk0J9gq3UwfbXMlbqc+Vod0hu2mzRFbdTWImK
ipM7NcJvKkZK3Ni6a/yR2LDGZbzEnjKwem80wFjCxZj51BsKHEY5LErc9hoAd535bKHREKlou14B
j7+ZDAAKcXEfJjfLYT7xu14iVQGO6X+7tSQFWPqDyTKk9P7hNHP7GsQwGu0DI0did5uiZMAcGHlR
ku4ryDahksRTVDAoYFaRcUbfkBTgT1zhrDGGR55srut4RkenMmqWYYDjKwaGLCb5xbLlOX90GxpQ
vSvhrV71NUfh0FSuuQiJKMUqO6V4FObYGK1IDVEi1OJPoY9/C6UQOBJwNsg9Z6JtOXh13H2lEovS
lWGDTfTb9yj8RB+DDFpZDjlAHxSkd4NBPTBMFv5iIFS3FpMGG1Pz0k6f7urYW9OMsGPKxeyt/xXO
P8SPhGug3VMmCXvoeziYL33I33scljk/xzKHV+y4HLsmLAgHHp7mmQOFUf0jQTP9phgiP9Kh87s9
OXsvEg5rL8jYZ49KHjfQdunFm2TSI8Q6HXAVvKakoE7DYPo4SMQJLsOuJShSCpcoPsk2p3oUbp2l
TV9liM2SubPZz5GgTNM3uzSHIiV/U4jfuU8UD3HJ7cdxAvEpbsDe/ZSlvMtxgYlevCvw7EAeGQpe
7WKymHAXIsMlOEk0eShMJWL+lMQnJEUobY1QwYLSAgrXDrYkgjrKlREBjy3mpngwfh72rsLVwIKc
JkRNNK396w/Rp8vHUyftp92qCzKp0e6VYw8rJm/PQvehXVWtiEZt3+Bx8uz//LVDv/5EvXF7VO2J
Yxp+/9By/lwsK6thvPgyqS2czTMtw64k4V9b6O3Bqd2QaRKnO/+nHMfKXasO8622jIvltDY9pjja
adyEQUaHICwqsqp5UDh4+L8lXFXIlWuASE7LpEZrlnCWkzKLFFdw1N0SEJ1stODqf2nTN3z8Icx+
BQLL96lRCthl1IcNUaTdDa2sL0MRARGI+IU3j6AMN7IuLbRQIgfbojtH4jlgBlnyfNLWCjQlYrvB
ZdEWnnbNk7Icr3XmxIdtug66Zt/0BcD/orzsBZ1lXNtroDdr4JyrCEfj20KPPFlPPhbplVNPMCbY
sOqejNqVawPkKwx0okBK6AAZ8BRiAxdlvHsSGXEumekkFj6JR0s8W8DDqBNHN2oVrlhtdAR7bsdl
lIPAxHZ8REQrNWli0BR3Y7D32EAR46NtbJU95GQYTbylXbkS87sZIjeaiWLmhg4bBZ65CPqOa7hc
1z92nrh2aeGQCbQxXu2O2bMrtgBuafSeLJd/93wPGqXcXsyUEFvIR+sLOxF+8P8wG0jK7fDUXLnt
qR9iFofrz87ZixUV2yLu5yhtNwfiWlNKJWwhuf9w8lEVVZw64BLfupi0eXHXDTt4CBEeOpD07CE9
M9Re5T+ZybpYklFcJgSlpD0GFlvcewgimZUJsp/G6uHoTXGwY5uMX5/IP3vTTQLNqPbaPw6ywaGP
+Fo0J1u1Z7HZX+CCNZofQVrqUwOJQKufynl+syCXzt+gXODIsjL6ADePF4F0wsWWjwYV4RuWWyaN
vT0/Yk/XGQVaS+kfuJDUs8Q7sIcaW6ZaiD7olM2iPonDJ3zheCbkM3A+A8kGZOuuy/oRzLRYidPM
OHBrTVTkh0ndbQYvdlQAE7upufKisfQxgPW7wOkxDNXvLUqAcmOd0REwblGJTmZivWYPLAcc49nt
rEekllQQA7K8myNPZoo0bRhGgTrF6On1fW+8RgZNhI6rXy/TxODR9bGa+ckQbfffxNvs7A3xTsbw
HsPpuSa0i8I5St+AYdlwoYN0BtHWfSVzRz2PIfMhgXrPlD2HHBqYNUfbQqkSQJAfI02qXhK9ntTz
KsofZCwM/ke8ZkEEJoCMeMdU+1Ckwv8bE8hAPuEKNbAFf/YPJ2rgaesUsdU7RIlRqwsx0nk9B0B3
Rr9mv5BfYtXkzSjR+N+xoYQ+FDv9lvI108bufx1aUEZfprwSH1ZG1tklI2D2vAvMJ9dDq+6mQqDk
kTCc4Jaeoyp/IYrahEDD3hyowcN+EQiPMt/r95qGmcJw1aFvmpcBhQxrWYYu4ZVUa4e+Djt9+9P1
hy5WkcMR4k0c5jaBz79xoJR2xUK+pTD/SbeFQRU8i+FSh8j8TxWMsgaclTk7jpWFOg250ZjXMGhD
E11vn8ZATcmVXXJqSTBBIqwqiMya6pls0ImRcT3Xr4/W+GenSYkkqZEtJcq1tcSZ4Sjb3iiaMXxr
VcM6aCQ5eskW10QxBOCrFIvOpaV+A/aN1Su2znvK7KjKf7uS6fg3inAciShrmjxDDUA90KXSiURu
js6iDf6qAZckgLJ/qxChmPFD1OmohZlss0SZEHhF7oZcdIilhwrciHIoC8Rm5EXPp/0PXS0wj0a1
UZ/or/es0fExhvCBQ50SVITjcHvnOliS1kE8/VkqI4vKatbOj7qguSW7d7F4trLMraBonSeOyPW/
HGQ5XIFB1RSGhQ1KeGkxfo1EAze8M6Nj6wrSDT+cEvTx8QsSgdTZuty05mO3jHlxqR1pnmkOu1BP
MxnhD34iHKcbFPpPCAN3sCAkR9WHjX1R8bhg5jHVxLl3HMvcwH3nBCBb8VcTC+pVuHIOGwVB82eR
o8oMKoCQNbS4QyhTxtQQ3eODm761ylP4Qrqm8S6umVEZLYp1peOvETy0S94BTj3+X94jGS8vqlBD
7C5PWfg0NlVihbD51mBhi7WcVUATvP9N/gdoapo4BmtIXPNVOe1IhCD4lOCDmDZTIv1r6FPjEAfC
VUBnUwSILfx5lNUt0/5JCbvd1JKVhsvAhyic6VwP5FXJgNYO56jAAnpbnhlzHDLJstXMbLKHPwt0
XoDz8ITNLhUXJ/Go4ev4i7akAhDdOI0SRSFd8X2vkh4sES0dn4I3n9yy1lWd5KtOCIIgek1+n0qD
Kzrrgbn09jO3nmw1j1kKIKrd7Wi8lzCRhR41YpxtsAp0O8hCZwD9bFX3tZ7NeNMV7I25wTvVGix4
ykScoyLyCpfYFAE+2udK0Jo6dtJuYP7jtLhx5md9Rc1pQshsM0KLh9EumFAZXtkn9NwwWwoyVbiN
VijNcx3gG7+C/KyzhF7ybela9iotPS+Ff9COjOOdUCP0ys+W9DlZiXN26QjUKQiSkNcl+JuELC/H
wSGuNvhjzOZGPCSU2UyGSsSGdyW2aoHpVVoX+Iu/UhHbGgycHK8LX0xsHwIoFoM9jNRKV1/d/GAv
AKGJT251IqV3eFhXEZ97dBv1/B0OyVn2lU7khlmiMNUCePrKn6qEKOM9xJ2eozoQJNQHder+FABz
2mthYkHrqGrHY2F3fpGBi0wgOEwrS5ExHoyX4Mfr8rqAAdunhC6TEan7yeHWNz84f8ZJX3IKd+gQ
whnaLH/Vo/agmECCJfCl41cj9OmpFbCVAzCqdo6lqHcD/yFKaah1bErZhRRkaKCPa5+nInrIt3ej
SL8gFj6bJhz378DflTXVzlDWw02dwy345Bpmr1AIfwhWm9/RXP+OTzAh6mX1ndsrOvu99uM7wozc
zfKJ2ly5wZ7mrVApQu25XwkOGayrnlQQaP/ZIQOozIyVfDm8kggWl23x5t+DzninDEmg81uvRfWJ
zuuwTlyXyOoKwZS4PgKSCzCMg3l4RhahbBlZBzWA1CWjLx4nReIzQJ/DoeLNzn620G0tYHzTCnr0
mipc35od/mMOxqxfSH9LO/2dRfPrnZN8hUVCpXejQlzTX1+5hCo+cPwVipsaZFbaBzRcTaZPvnOk
J5now00k+lbXqPPf0yLdbpDkxoDVXL58BRXsk5PfmcJ8rbRW5webu+dTW36yk0SljfQnDAULKlET
DeWeUbYwkE6kHLl89p9pzV/URcOUE5fBOxMtCzTgl6UdZJTaq43fWRgNRnQw2K/eDhdiC3+YyljS
1V+k0k/ZtLUt6ypW8L2v2fkEojNUZJDkxdsB81fleWtB7sXafoTjWfnpEfm8h+G+JMQLWHoaKB0B
ONbSCV5Odvw9qxW+fCrwXvCoJCI8DF1oEGpkh8pobSo6cwlVk7H2x73F4sGZxvWR4jVBy4ubL/kh
HrzQV4PoQK2pXJrfaGKyHCu3paeArvovhRJYLDC2gIs/NLECtisyA5kkKcB0lmSYtWkyuIxJQBpM
NmeICzYLqKVFoo/VUgqow6bXxw6DpNFgV1KAUgED2BwZqip2fRUnrxnVpDa2j1cPzGOInsfALQRK
0N+G4aJRhRA85rOwBMU0KBahA2ek62u+E6XOSRwaAhxAom3fD7nbSZwGCi1Q/zGvAC1OVT6fuZT3
8NGeQ2vMbuJnieDh5B27xNB4mphA+rMFTXiCXwVvZXoCZlhyp9DjPr4u9t9zp1/9PwaJJYfPvuC5
eMMU79VoE59jx95uGw9zJytcf6/aLGK20NCJ0FwgLnfTqTLNM4nel8wRZXAjAYhFGnIby9m9dafk
Q8QNAHuxxo5Kw4LY6ApP69x3VcY8JA/ag9mGU4xjqQml4fH6uAj7oKd6qoLfPtns+9fsADl4WJyk
NqIUvBop+HWTnX1ttXIZFN9jg1QGbmUpKF/OD1qaTxEeDvgFfvsrxKcUOm0fgylz3tsErzMdQL1V
s9I99cNz2tDtCKiQGikG6Jb2xyQODwxAzOTBG8FVlGTATTdJG0uZzMOJ46nz6Fm1mNS3Rx/lQMGD
V0c/sh87Wt0W6ayx3rgYZ+hKn9++gJ4vr3qYc0jDQjcwSLAYDykOLWZzyrs6DVr5iBLSG0F5joGy
dTSfzW88zJBFNg93p98bDwd6VBrM66D3YftLG+cFPDa8IpjBijWdukfYUnBAfaMcsvZOsuvfhxbf
jd6vi9rftW5lyVaRdbix2cprEOJPzBB0FD7QV2vX9KdZvqAjs+cSURXFWVeXtx7wYcjYKADiMCoA
+9+nnc8zucHD/wJP6VU5LENfJdf+K3hG/TlBqP0vpyB9hD/S7wcDSDMrA8XobOFxKJrW8VCYnkOg
K4sBMe0K6xns4chsyVtujbIcB3TRJYdk51qOhf6pOpF7Tby9zt95l4oFQsSu0S6ImMmdaOPscO87
t6QQTiGdNIpmbtrxSlB8uOATi0gwrrJgSX9R7XmfblF0Iz9GtlW3tG9psOir4Jxm6xYqfvKKdZZ+
cuExYmcoPNx+fYFU/73lonwKfRtaE9j0BIaS3EXa9dZenEsfkydu+ppQ1euRVoAok2XCCafZiwA/
e6hWaLs25vNGLsfnZkH2ohdc3NsE2PTwQDjE3RyIHUz4klEIPfIylr3zw6pIGo9PozLKgJQjCv1M
rDVjespj1F1qWrR+R0eYTE9GfsE6IJDLbcEuXC5LckUwuwu6x7gcgzDHZIpCrT5c+5zxksZXmmmP
h7z4iwo/zHiUS9HHsr67l8HV6zItyhGiflBakp2QFcnYxPk/ZyNV+0fgjUNv8pTpOmGdsXhOMH0R
2lEGDffhEXr96cMlcdOQz+0Zkr5O6oPbHxJNQbBGeYJtnXxY/pYBdnkGyphaHxr3wQDVGhnqMLhA
j0o4JzKKOZl2GOVZQTvLQUE4RbTKGyABU54zGxC9BHXpELdUXwFxFOsNVPbpVNwUS1SKjzflwI51
zSe6MrQ8I+PCpqCHewsByiSA7TDbWUL1mKhSEhl35C8C3LCqUepmc4OzbIUZRjRBxMy+ufbuBFVW
+c1nAqHP6J830PgwR7PWo2GPlSZ5DkcXgiIAgJdm+cfCU1nO8YLDkI+tn6TQ7+2VS6Gg5rHCbH80
TQNkKmk+GCfVGg5qFFoDiJrIRh8Jq5NwLd5LPrWl19LoBMSQzn61dyfviaVd/GttzUUiLUe71HAw
tgGpyqoIYo6FIfd3uit9a89VYOW/gCByE1uEkvuKbzV7ZhKH21X4keH2qi95XHakGPr1mSbcr2VX
Oxa7x/8rhVMTAa03Micu+xzGox84mATY6dDjo4SZ3NA4xkgKASiNvH4ftKX1n2TD0ODvFGCQNEu2
gCfWJVCJ0Aj86Wi5Ugx5Yo2y5Y8kmDdPaXZhc0cTAslS0mkYckIzr6JtUNtrhnj48Vxa/GSpUR1j
4UYxfVhhfLuaHk9F09K/8mUmuHF8qHZ/ShUhn3QjVEzrCfPMIGKkePJ3Zw0QQk42xNu3GOJ3Cxrb
0BzgKvQLLtO1kGDYQkmML07/JJ6IL4CqCNEu7NDzd7OdOa92dYW2JLgkDJojuVQfGf7epRPbR2aI
9JK72PERegtfGujUqbFDKXTe9znwfKCUfi6WpWWkFdnRDv1AidPZe8OwyPSZmXip6DyY5SZd4qwb
9HjiTBaVAvgTcf8mMb+r3CG5ktCSy7gZ7i8GTQ5TFRE7aWTsVV7x8SH8C1BFc7mggAG6N7vCIRds
m4gDMo/SClgF+LGYY9i25LG5wC5KA1w=
`pragma protect end_protected

