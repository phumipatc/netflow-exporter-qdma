`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
aV4vCdvimmJHW1Ue7QMkcCc7SnRoBHU0aItImDcV6uk8Y9iOT8ru+mLRRCr3OURtyF14o89WhFgl
kCSwEo/IBey0c90VF7b/eWWXh6l3+qR1H7OY8XxAwIss60j8DUxS4BZ05bewT7nSBscmzZbuj5FD
hev7sUOt64n2LqJSr4b6xkFQ+Z+zalgb2dpoCyqx9CoFQ/hoVrzcEn9J7cztPfcqcSn5Vo81meSh
Ty700KQOAka3oNJMC9PPRZ3a7h4hH4nJO0DRN32WGIAyrs5t9yxkmvZz5D17MOJFhLkeBOF3rreM
DdCuZj9t6mZ7x8Q6YUgJUIhjHfLmZsqR2D9/Fg==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
FRDGjAWDGCV7ofnnb1Nnu9gyLC1yzdvWSld2o0aucEq1Ku6NvJOtWRhXxFFmLPgowokXJISce6tg
uiN1r2FcXKVLD6rpNfTt/zW59u1tdvNukb0fSALpJN0jJRFQealkxzQST0S8+o4uG6IF237HDtDN
ieDKbCQ6rqu05jZjQEQLic24YRGljBzwgwwZrt6sq1+Yk/SY9U53yjze4rLeCfgwyyR7af6780yS
QsdvDnIfkOBEK+MfkW7La6EbjEtOWvy8ueGx0g6oZdvkY8tMKrd0ZwhAXWx+oqqqq9lQicO/jOQQ
GBGEhLd6uQ9+DQyC84CDYQEmxtMaMv0n1VYP5wAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
VD9l733JPE8sGtU2SPPQGq5jfSgvUF8iOW6yjYGmRmM71zsUor/7I1TiBThCO4yrROkQuuLRNWT9
QscoMDqRpg==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Aq6NN8SBacb06NEeh2TwLXfydh/xQAeuV1/sTArj7NlcpR+uBaPZ1vxQFuEIYjsxIcauh/yJl1bn
yTGo6BTKCIUYb/A1h8/KYENXQLmQNCM+EGCNa9aOIetbWp7xrAB0e/jPLLMWQZBBET9FMsrdCvuJ
03q+6BbOjFphLzjPvoj6HbgAKZaLXKpybjv9m/Ar0TueA5QwmdaFZeG6///CqKzt0etEG+81cf6j
aH6wNbTnrA9CMX+FpH70rbKUZYHDVBe1l1IyDUvLuvbAIZGnX114pMLWvC3/3AAc4ARApfM5zxCy
GHh4fhk/y14x8yq3P/3tQ5J7UNUOnOHEPvy8JA==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
M61BQDGKq5aE73o8hlqn8ixVSmKfoQywscztFBjBHta8wdSyVkq3okOI8vnjLYh8cSkc7w7/VCu9
Jm/Kotfn4P5L9ZvLIu/8QG6hsv46hUhycBsb73ZhbJz96I6nuTM0HLwos+ctfwBNAe3tCcPKsALt
uwkbM1ghzbaPIdjDgo2WXVAE2NumIto9bCx9kZsnE3iCNLo5V/wpkJpStACfUowNzG7agRllxtkk
KEzCwuzo03K1V3Z/uyu51CqUu7ZQZeEzdhwRJ+XACQm2VKBR1z8IrV4qwgTPhkHymCy857K9DrAP
o9BC1zMNa0wT5VXS9xCm3txjivPNdekdOWFx2w==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
WYKtJDkT/jCP7QQAb8quCVydeZCvAdRp8/cSjkuH+8Xg99ORh6UHOaJLfqDDkLOjCGQ+SnW4T7+L
SQ764t/NcQzWmuX0PhWp3O26YvKniyTTxFe8OAW4MwXnd8iYOJZxPg0ObdzHgmZKWQDckG02W8k/
qBe9P+tuomSQijIxKP0=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
p+ns4nzmPlHC0BjSfOzJA9xxDqNXcjEpnYoNv/JtJbLOdbf4tphJgk3qcEl4XaHCWkkVguJVBt2Y
ofB0FCpEe7CCfLgKGzE0cThhIX4N9cKgqe497z1Mr00hDkmN4YDEKgm2ORCXc6U3QBpoP6JA5HJE
Mj/kfCMA0pHsooMyd6DkWqI6WjKFJNUn5Qf4e5u6k6wFNKfluTU8AaAfPeRnENE6FmJTisIMMXO8
5I7UyBLidTmugbLJoEZk+kSMkpvQEJUPyKieWX3IJdlwkIaxs2SRJLc4joV7LP0aImq7MwECtdrt
br5UPFfQQYEKXol3tHjrwjMDVdbRN95lJdPaTA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
2zTfrqAeEC+oxdRZJYJj4UlilqlJ81jq/TlKW5kU75RKBlKCN39pNGI94L7ijCYGmijdGXxx1Jqj
EKaDuLRzk2XXheOSPwV85oCoAKxFHPAu9N1XHLpxWkwwBmw3gfyeoJPC5+mDI01+E4HHByP9TG96
CarHMpcjcmXJT7svqQ//gbs+ABNCNieqNM1N2bF8fnC1l39ywRorCL2bRUiyoROQJk5VYZrajyst
uuX24HFyOxzuZtk0i2zDflqLxlmCRl9VWvuvg5L3aqz0E2MWksFbogVXbEP9VE+IKI+S59n2Bx+H
VdL61ThTeI+K8iN8SRqCiT/nOeLh2vKu1x69lQ==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GHBuBMpwbocgwT3sX9tC1SrZqXwjWRWI//a2eUGfSRH6il8FO2LVmHSgOqU+cm8UrUmYpBXazHz+
7dzDRPYB+OX480FIwwIFopVeasoZhnd4QjGzFAteM7ZyTU1yaXNbycS66OPdp90LdbRsYkww4z1t
tH+g98eZ1NpEPLzCDbE=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
fymI3oNJOy7NXtJ3Uj8kVaGkcq2n2jNSWWM2VhpQyHlN4aiGWJQfkOiY+hIg1ZRtY0Psgwr4o+oW
5ZHkpkm/I1jfKiUlitUifHLJYzpIJd2M4/VohRcFdka/G/4kJaxxQ4q2SFtNuWQswCHT2zyEQ4hx
v4th0vJIK2WJGspid5FkN/x9EMDEDCleKOlKddRWxrAOLyd8au/WlQB1kOL90iv+WbiVS0rIJtJI
EpyHcR8iZm1PAA5lbowc2HRJBnCzSZ8ZoW6bI1rOGHfbw3z8tZh8HVUpqpCjVs6gAQIuftrD7NhN
lukWQBS/cY/NVyFSr2wy1Mq6NHOJYLru88hkUg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 32288)
`pragma protect data_block
kpgXnglEvbZefDSoRBMf26i/eqVvHvxZPUsIwYdimBYlznI3A4q2VQeyCtagZfjYK7Pt/LzHNxUx
98HXogItapnehnLh3jN4601RxEmot0ziNSbv4z64hc1AunIRWyyHigYCs4XDQkYVvNlRcgzi5zcs
1lOhHVJfEnd1qv0NE54T2eqLixeMYPTcS3DusM9+ko0KIPEMpxctTNrl7wqzajwVU5qw1HQGQiuj
JUkoHjCSn2uwlmo5ojAtRAr+w170Dp+dgpoWQTl3iUawUrUdqHyfxhs0atRydocVHK3K5ezsjNO5
ikSd64KZ5GsIdJfgImr93L9hmZV0CjUbf2d47JNQGjr2mX6BLcuJTkX/ba/CBMzdrF8OFRxl+giI
YpcVTL/jou+Wp+MOQr5eEUmBeG+OoTojywxuezhPPTB+cHC0Dv1M1abr5lYIAzAtKuHGm9Osu9Yq
tZ0WAVFtSeLFOstMoRMRu91SV5Z3vw/JGuwqyNRNDG1+4ymG9pnHRr2RJ2dInx5rit6jNYwRLl5+
46H+76DzHcKEjKH5AHCu8EbaeypVod3yedVEfqy4FDnm5E1N7Ajrhsb4TtOjMtbU12Nc/GuCHnfL
QkTr/EcuhODobp3KuLkNiAQi57wclfawXXcok6CVGV6jIA//Xm+0JZOsoG+Br4/V77skeBUNHxO3
jDYsDR8hgRLVivpp500uNXYynGz98UpBpZ7I+B5jkOnpFZBuQxZvGf2JuSYKu7U5EfQdzmmyIfyf
r5oOpgQP1s4yvVx/B8WwNDa0jPUTYls4drQHMy61o2YPro8084TRRo/lzcRrPkNS1hE9Jl/F6QXx
9/V7rnhVQARqJ6YrMrEKwAsGkK5XpIREdY/dlxy6pCAv9M3oWvCt7UoQ/hIV/3nz1el3L4QDmqS5
irVbwNhODVDUEvGM0RcpawDEHKMoxam1HWom7lEiOswqP9YxOaVSDK3ZpmIPZQ6SPUKQgWU3nGQu
eV22bTjrlovo8sn49cJjDxmu423un4kCKK5TiP4z9yV8ZP46bPBWmhHxaF5aEsCaNdsGS8ufgWq3
NeKGV2dXgQZ9Gbo7oKZXw74IjWa4KnT739SnLS4VsJ6XDd9xNej8m4nwkZCNwytJBNvf/73jZSkq
ss4/ImFsOdCzuT8rpXSHXt0xkm1MXtqjlNcvON8VDhxTAT17Xl1AwyiKm7CgB01vmLtMl74EbG0X
8aIayN4gAEIvLGIeYs7Qeh4mneeAlPq5LgNI+DqrYqVfG6iWc5Ph+07+wM26XklFKOOAEHiDxwBo
Iyi9l7cHhNfuF3R1E399vWb0sq43QcRrm5yIIklYddy3CvMKxtwnJobEX/LVB2zjqeCQGkodIhFM
RomgAml36rqnGP3c4nq+LqYXqiqiTd5ah+iLHgjcR8TFm4jbfJQUYorhlKd3OLitGlU89qlwPtiG
MNiepWpB5/jhkuN3By4hvmI+OYimVndgAP+vndO0bRj7y8/VokVbNEUlAAN5WH0L5wu9BsPfFO9+
hxz24GYfgTcTy81Zfbefqkh9BCe8M4CaGxzTXGrlVV6+kl8+6DlaXdsZhJkYspnWBCtr+dOETI2I
wxL2HCKbKy4jPPNycZ0pnzPfooybbqwYxQvB9keRSxej8JUgEW1m31ve9E2ga5NwZ5Q+0Zor6B5P
QcBA+AcTEZSJJjhZoEVlcURzqcqCm3qGL3iMl1s2UDyw9cgBtNwuiI/fKFo5GiaB3l5lADjuvmGH
9O5oGFsNPnNN8T6+wUQ9qanPdIU0Ecy0qnLkYY3f4jxmo4ST8w0rNecKdJsRQART0p1Q3jCIjN8S
hEIIXxDFtdKj5gW1Mgf2HoTn7LjiqduRwFhmNrxDsXR1+K9GgfpChZX28gHvS/Asm1ELfgFTr682
VZATe+vX96bfxpk6kw/kUYcHUwKtnl1EXI7wBhc4ol1piO9eswAaupR3wAZnCmXKbm0PG7zxQbJw
UdTSx1C63bG5OMziPjqoJpUu8r3B1EakdhkMT7V23ihpRv4WDdRlxQ+Xd5wx7lAJNsyli9m9JLgk
IAf5PHqD030eE5V1FnY8yX9Am7QBJXLXA5Aoznmk52SapObg+yO8h5jZ/GY3LHImZJVyXzKNIgM5
hZ5zTLYyqDmGUtbLX1v9SfDPylzJG+xwzVTMpkKfnLfp1MGBYzi+X/kKTjw7FA9Qj1qBd+G74z3t
4L3k7h+KC9JuQ3iPnBaXm83sg5e2nJ0g5ecNWkSMV1P0Sah39FZ9BPfnGxXDOMxOQwBHSlyAnY6g
MuyTJozKFIcIMT3WeKROvOF6o08xweInCNyfYv2FLdagWzWMYV7ZQs2gAKfA4vhHbUvrIOU0Tpwt
9OwMzgXYNap79PV2GtqqyleoQJyl0AZwmYODmG79pXns8TxCTfqk7CM77oXYkR/ZjY1ek55sNqhw
k0SF9lAMY6Fp7bGKBh4kz0PyAeQggouMb/PmViylvU3sRCuKCeFHcwJmswV/1l5POQ6Brb44erXa
2tr4eYsAzjVr8TDNqqt1xzkm9UVOWhLiPPIIyud6MAb849VraY3qB9FaLxDT/irdBE1Xm8A/yClO
heceSZvc4FJltoX+7sKxP1RSoWU4agBW8rHpW31XH/1r5/uXk0yESAmLutoI3U/VLV7LlP6Z+9gp
nEEwwEDM2YDxjoNzAXI8omRCrmXeFp7nPTPjNJdNOTdnRDUzEvECdv7u7+fj4RA5kdAwts6itzQi
I5DMu1p08di8KkFeBczTpyy8hTHUAvnoaZRF9LCigUfsAxGjeikv56JC6Vr19d8ALlwbVzdukrjp
8VhPc075AClZx5GnhDsdecamYNSuh1AnrUh+2D05BgbX9w9h9j7+DfJHF9E9RApmlzM4KqLS60KS
H4H0tVIHkMulRiVyit1Vou0zkkr0tjztkvsbuhvf+Ep8xU3CJcRzkI38d55r81/N06s/aT1szMkD
NhIhUUMHwMxAUVm4njhyiJCb/5K7Uac8bq2USoMGBVlvoceacJgZKmj/H2SxXA5MwAmaZGoXOm1Q
YyBUSQp3Ec3SBDkiC4aIC7WA9t14IdRZ4salOTJrr7StB09tKIDH38MMNJYZc+TgMQpMaIxhObYO
wnXG2JSEdY+hM+Dpob/OeRvn2n3aSiuWd146zV+KBIeAS83HkbUtH8eLfMS5h1zUBjiRyKcsVK4u
6CO3UaHw3iF0j0RXNDTUNSBl5UlAIXr/8qv4TIucjvxKL7UW+oJsi0Y9AN9DIzYy9UgMfM48Oc7i
7lqRFkgGnaDvKnsIuRLJDZlf3UK/HqSTejFlll8R+znHQbT8dzpEwUqD99McAbXKUOaKVk619Th2
s20fNENm1jxbBOq/aj1JCaoBMQvEbTV3aDoavhoNWUzo95E8iv3XH6T3vwO17vezas4cVNOUyGxw
kKK0VH6ZXS6YNQV19l9spXD1vDJ2RbhzXLHJAK6+fm3dtwsKVwv/dMxLEgn+X+5lEkiP+Salbbll
xv1yePsS37VswPOsqxalTdDZhOKHuyTEt7I9/WDg1CKhgUyCCS7azZmESj5A5CQ7mbSRrzgprQf8
LIFnctObYxf37v3MZEChaRrJA82nXKlcryt8mmQtNfbNDtdeKBJxdVHWE/lXeoH62zULPm9W6Krp
s6yS6klFRLKF6gMEWOJ0KFxCgg9iRZASoJ8wIxD5+Y01vSvi8ZERwOQTAKd6jBH4e+jWMvs5pDnE
wVRJwh7hOHUJMDqeUvX5aYvgdV0HKaqwtjB3y3+QzyT/eRggFULfcxlfgui47SutUBUgp4UYOAZY
7pve/qD+BJ4B0jqTmEAbI1qjRkHIM3DNa/OmZB2pEVRaW35pRUoye5KQfRo18jOhs1Ho0Ea6Wuim
9+EZCiks0qAFMIje/JXJmIR1mwv93T2de+DKbEE023TU4MDNmXFPqjmipqkP9j7Er5LhV1q5meax
xy7oamhGe6xVmAd5xIKBEiDgWu5iv8n8was+iIy6O+G7iKukriowGa9Rh6/yF8eIbhuyDtQ42bD0
gYKz5Wt3c8Wft+zlRCjgtTSGofLpf2fbQxY0EfvkZ9falUkGFIlYF9TPbx3Jv5SLXrlUbgshc4UF
GkqtFgbwMSm2DuhtNMvFAJy6oiMRlhwHn/jZXdmN55vvLxE51GRyBcnvMzq+UByJDPSADTDChO2o
l7YttqJaZS4YvIYRNGaAg77mZaAP63/F7r0Ve59hVKZQZJBx6cjXXvQrCB7i3FDDDZzIr/6Lmuar
ZHI3C4kXLBOgHUFwXg+n7Gy+OqoVPKV5oHWr+qa2FzwEmbbEFVefFeemFFbZXQgiVmy8QqZMpsOW
ysN1B6BNRoEatkkJWYCAAWoVSXzU0IyDuA8MKs98wC3woqnfzohrJgx/9mI5VjbUn1Y4cb1CVZRG
rlOmC3nxIDeoQAELiv1Eo/qs5tKGQGGOg+HvWnEjQw0NmrxbRTkqWx8Ob3FcBEX5ESTbtg3p4uUG
FTZ+xuegMyKvpOfsfcip+77Z440JirCCEZaja8WvyDZJpQc5/0m9L/FzH3bCYi916jk4DprR2108
FVbVBsScTYzbyczuslhFWMYA8dFNC7Cdv4dPGh3B9LB7cj1z4GlUwl6YcXZsjGRBNb6s6YPEmiVX
lOb2sxTVlJyYwp1+QR9clGkWnWrxys5U8sWgizV2Tao2GASa3mv5dvy+FbCSEo80/Ap8TckDojh5
POIt8d8GVDIU7ZXokKo0bYI9itt0wW5uRxQMtfZJ8uf/JCuSprus+j4LeTBB3ud225rR5TR5ZKIw
AmLj4Iy+mJTuPY4xS/a5JCPp/ID+pQnYWTwk9GzuOzwCeLRF7DrsogvTyGE8igag+RUF8222AvIz
341C7knJhQD+x+MsuO81fNI1xu5yuDVLG457JnVLDwhtGGtj6DCBgVILe6wveo/jnFywM6hMQuWt
2unHmzT8UI2SUou484bKQ3oz9ykZZjjpzY2iSYgY1mlfiw3apcj/ZjmhA5GsOYETyxjRsFINnbQG
2s89S+Rt1VS91/Y/eOS5bVI6fEfRJPjWy9y49K+IYR7QzUrsxOGoV01aoFiA9F9r7rVpDcsqRBG1
89K60bIlJtoDeTukUHzmrF4ilumiVKj1RGb/ZKoRfR1K1qUwj2quT1teFNrYOtL5Kp31pVN4+dhB
oc2JPARhJtOVNMCLo1T/Wle+bY9DdMGetHeDQ+vBI/sfeCbC3xw4mEwEGtSyexsWsIOXcX4FSdgA
M7TPm32z2vlFvDs0rcRVS0jerELw1iCNcNrmM9t7wmjDUaPeXTDF7Pn6JIrw/7a/OzdY4NNQz9Sg
GmHaaG7pp91Gcr+dl2BULJaFJDH58gjwUcjIfA8Qt86VCdOHQ9UxKtjx6bMnKjSNyiwXbBGBdj4Z
HnjzJ/HQVoyTYc3onuI7H1z+2hs7At5sxur5ccAHnD7EUSWRrF45b45f6elHHfkFbYOHIIszCP8E
pX4BVje+gKGRAEFhLORfCiuHK+J4dBnga7Akl8Uh1MaFPFXMRqgvvVNxECAUEU6FfmqnrElLEnga
jpOUJstNv0S3srWw7W6XsxL/C8gCQ2IsWJOEjsHa3ACTVu8y4J9UELg1XhOSnOILvnAUahvZ5eoC
qeYPeK829LQtt9o8XmyQhkdwfbCds0VoRi9cpJhg0rfqr153gFftHClHLrLv0pWHtkXy6YfN4MHY
4s4oxpLaDH3iu6Sxa0iqqs/WdSOtROmtJ0rRfVBAkg8UT3r33bSJn9/5689L4R7M1LH4I9wuCJAx
rpJCKAh9Mh8V1zG+YOIyWuZSUz9iAZqkIaHpEX1YjA4BDN3UyuaQtxOcKsFVrHs9dN4eGLpkLctP
xBLQH3yGSiTEuzp095Fk0FS2AACYHUd3Wr/sO76OI9NJ8LX6TLDDm7WD9WU7kjqNrlraTcPaRwJu
iCaXwdg7CsyCmFfVZWvpAEfPy6Df0gARcs7E2VTkaFzZHiU7NBW7bgP2D7QsEs5+DP6gfdNs2fod
FJiWI5J6hT3fGt1pzAzXky9AA5tUP8B8Pa5nAv4eSyc1MuHW7dHvk5QA3T7EYQlzITnuReXQxMaV
wdarbcrb96iBcqw40jHvSb5hdlBw4XDbphdGB48+stkcE+hhDf/n7gid0SSSPHLuKBSIGkOMciQU
KedpUgrVvjmSuCk3A5T1rz4FMkL1XbLuaz6KTcXnltSsEIK6xKb9pHB2Na7KSqXu18uamsb4OTCO
oka+Z5ZoTQSBkqIVAXda7UZd//V/EU9w9On7h7DvSa9kITxHHPBSaAUGqlATw0+XyTlnWZqQwaFY
lLgpQaEN43B63Nl/mK7fOiNDg7brtOl/nnibRDi/2KZrAr0RB8IV3yPBUibiXW3YEjE0jZLxcm03
UM0WUvbn5wKGm95I1yMUJbYlctq3SCF9TRoP4lkJEAlL7dafGT5QoFOv+nuo1prlV8wFdPCJ+zQ7
O1eKzhF0m+zPfqjfvKyaWuLXvke1A/QRKcKI7PQbEAQRUjPriFxKobIkGxlbF/x2DCVZTn4k5EO9
250rneDHpBwDFd9WzYlxVWCUBmtSoZD9pF21s0s1svdrWHi9P54LIEcwq64cFVuFC4sAIqylja8z
XZ4coM35lXq4MY8SofqS404vmfi3Y7LgQcZ3zSSvsZazqqZILFUxIJJDlrV6MUec61mFPDucvlj6
lc2KVXTEe74Q7a1XF+qIK83Dd/PFMfBS7XU7CsKANNgqDJ/n075+chM597BcHThqODWqnC5B/hf7
qxLwvEWLVU7IcgZFMsN6fFU/QE9TFoDEJDD41DPgus1oYm6xUHP0IdiPeUsKLAnr7GT/lrlCgNNB
8Zq7bZ/g0vOHdLOlWzslZJe9P+2PU/qDDTcwilcXduV0gKjsExJTNr7zgq7fV2kW33e1RL+yFn1/
uptliaSExT+g6ECxW9DyM9anym12xQdaXFbqCB6bPyI9qiIUbY/RYmUqj0PL4i8QvEAHum9mjmyG
/WQBUkpiiTQfXVyhlKczh2pB2G5WgQDStDxIqgwE+W41jKTZNxqUZHpmljraXTw1bn+1JTvT6203
bfuR9BID0o7RAsuqxkvyBnmuRhTgln6T4gp0B/3SamYux6f5OSlDu4ru1DZTeWhFAvWTCbN9S6+/
CRccqz5yZkr4k3sXQMl1uE0DUcbZX/rhSIrnBEJPuItosCFQ32f1WvAA64UVCwlcA9vomFcNt8RZ
ipnwRb34ltZ57fvO+yz9kloxN24SvNd3p6iiXQ2HFeNATmSczm/IYEuG/+KeqAFUHYECDGe0dtcG
kjc4RYdQcHRaZUJwl2gYbEJ96pok2K78IW/KIw+EFxGE5j0N+vTpZR7dDjB+brNwwFeeiKYW8gGe
W0NQm48QFjdrBGWjOAJlJGLcZZa2Hv9SkHlaCM2hTvxgDQaIoxNNDdu7vhcPWSrOZpEoRsx6BylA
VCHqhy7U8kCxZBszxq0kWG0zQfxGkKIC5Nx2b+59rTP4fYE6EjxERVatnvmbBVJwPOdw64iQlWAe
kMdzMlyeqdE13qgh+zQAzSSaGiWZ20YDVJSEJBHipiCrZJrPjDF53/6HV3iDjupc/9hUOyQ8Ru25
nzYYlGZZqqOkdPZ1PN9G57DdSetEue5jmRwdd5Cnn7lAv/cORcVOCIXlPABLhGbfxaY+7MTYRcCs
B5gbsNc05cDs2dW3Uwmc4TgDsQ/dyk0+/0hSDw6dbckWFV6Zn8HWKKsHBgcBmNZXjG6/S/jN3P+i
XOz+elBLCFrxKjdJ+S6R2TFhqQmtEuWWOl6NmhwSR4hoNu/gqeU40xISf+Iou8szK9rgcZLuazGL
b9sLLftxSQhL33qMl3OzRc0AnXWcwX0La/9Y6WBe97zkrqaUYIoBg1ZLZiBI2dcqBAZlP7V51EEN
Dav0LqqSaamAE0x7GCs9FmR8Xc6M8Dc9DB+bWbPliGsSgmXoeqe7X+xsm4bz8kDm/ytvfe/AOR+E
MagrcILs+Y/+cScfUwZgyuBeDuEKjAiD4XqKjI3ku1rlfvuRXaul4veLUGjmBhvdpEQork8vX3Qv
tWcfBgWLqSx83ax0M9HDSzyBK8goydFJUvAQKT0LJTuWDFPOtvBqYiMaDKVPt3yC44hjBqQO18Z2
LpitzjOL/Yik/vRw3TaALzGRhV3Qf57mIwpWrHJWr23LRSHv+WpP8CPfRt9Fs81jn/sP2G6byVVi
JOJTpIrbSi76GSVmlH2gTCFDG+8CrOaKlwkUmLyWvS9uXgryUw+OMb4ii4/foWMq/HoaMhkCqJGj
dBVGQ4WLe4pOXXWRh7Aoo5UvglmcOF9C8rBZviVedHXVAl7zsE7gwyj0/6lIJfPWf4DBt3Xqb+LM
aViQZtuRGds/RJ3nEUSHJzaE3fnD94BmI57nCU2K/Zye3NuomuUUZPX9vftLw3vvt604dmgcLKKB
fAs5aNQQJV3+tRWGrxC8mhvtggNAofUSb/bnm/jsfmwrU1LM6OtdBy6BgBahD8Lyq0biNNWiEau1
tRlBmoCRlHIV7IadmGNoZaAMpmYK2eTWJ0Xq6MiNISEs4C7Zu7OHvgnD9BBK2h6q81vmUCk5gNBK
vPzUcJ3j9khQ5nxA3Q/Rc9iVdozluHqv0bIzGg8gFcwDsvKwXbd90lxi8KBtsvdU68zDmkqKGOoX
2lTn69PR9jBCR1Ue4Tl4gY1RRL8/KZPQ1gcJCdwNWeY4H/11b/DV9FO+cCe11MOQyHqYWFXBjk+3
Jmov6Y8Nbx+hsUGblITfjaIaTb3gRbdouiT1gT5Bti0xaYGVzjyjz9GZSHu+s5VnP1HWXpottwwx
baCHJGnVa6bg0VXr+aC3BRxPY8GztBbFcletNSlz9HQfm2RVyXJrcoY5swk+QlsGaiP1yoWfdv5x
dAx/RXSwdbuNMPhFnKyDn9G396lzJae6p6pDrNI2ClkzjDxUULM2L7ZSouMFzAqHiH6jOfvbLLx0
fDY8xaj7HOuavTWetYn02wJUSvERGTT8dPOmvGwiLLtiRqDxy0GpeIkIFZHHXnMvtGLpjCeagINi
thwSyOwlSA3uLTf0ATVqpNcYt/4b1+bSgLOgyWlvmtERNpJItm6vreyjydjmuHxmh7ZZRlRqpfyj
hzdva3ooeeXLe9rFZ1rCJVtB+UaCNNDaqQFlryAiX+O8mMk3C+CzhLgxycEEH1Kobb7+nXNa413/
ElzVAQfJNTwcNzArduLKVSPXTcZUYNxH7TGLD4PasLgCjFHU3JhkVJIrlPclHF2zmE9qKfow0OqL
ET2prCmvO3ZdGx1vFb82YeuIHZpUPp85v6WdZJsV0snhVLgZl22Y3phkw2bazfkpFfOwznb7Uvx4
pnjg83GvzLu4jh6Gxg3HOQM5MQw7rRihnTIwSrX8x8Q5jvWizhDThMiI5TOvoJyWuxJ0reqAtAZN
h4NKEIehPmUB9lOxP10pB1db9EcGC59IWPm6VjNWmX4yTzAH2stODTHmG5Mebgr+DLKDftbDGIVE
qI3aqNKPLb/gdrwoIHCDPASQ24+QpStqeNEZJWBzXh4g9yXSw6u2TfKndO8LmBPp4t3M9mhrf6KA
UjiXNCl9NgXXGojRZ1OmBPq15TVhcCD8ntp3Prk3YXpJSHhFSM5PbdSSGTTJcDULadPbvnvpnrvj
xeEEm5J0nWGyTekqEhEzLnNsi1fzF4X8B9Ice5FXxbnE4WVBDPeQrUsa3qQJqUHfsDGhpxTlVOHR
TNAG6bK2se6IChvxU5cMfLcg+UQrMUlsYR0Qqp93LWpp93UpaPvx8WS6j3/jcjhp0YNqTX9O0jYy
gaDhwutnHnIUYXvH2Q+Y30M0clz23pkWjuizOIKm5HSm5G1aR+14TVNVg6znIn8TMKHTiidAKK3D
UV9B8KE3m4L/QJ4Dr6SJo0HlO+IOvhr7l+7CWFp67ZD3d2KdzrptR3JQFIIFglIKOzotoh0O23PD
UTPtTT9xIaf6sCEmS6KcZopJUqvUZRsgIP90ZorjBPwl4ZnPkj4E9UQ7EckOH7RuVFCXl+zOQgt4
s8vbDzkVO6z56iJS6rz8m1E2p5uolJPl/sOkm9HCsEf0r55OqX8nw0j3WERVNviBhRvjiphmJlGg
mGZ6g2Ceid2qQ6UAXkyphWBEw/a1a0ZoPe1WZZmNhBy10lkPyesiJHcXKXHkS24xyQhuvwcG8mf5
v4NFbdWJzYG+lnbs0GX3xUiPS+qUG+21jDrtLrFSlYJqGSxqAqqNpJQ48EvSmRU2LPI855WbFWDn
erkpp0auViVuww0kV/GqendReC5JCLwXGkzpO0e4YsM21JB8Cso8YK3ItdSyWinfrumVg6Ut91FL
9j2nMo5ngzIaY9HhDmQ3+glg4WBCEdP5mDlC7kRHAaFfwQxFVp1DQDZKbzgJ4sXyoPHqJN/Gwv8p
ZBwh+NdSzKm5qOXOlMVAn5KowfJi5/sqXr5Az4rTfRhnBMpD95q5rmYaNoSTKbARARYaPWVb3BpE
2dbTlJTfMeb8iRttIAnXj3T2iwykJiKSdsM6N0jGY5J7YadzCUl2xH/RC/FbFwCvHKTEem0/g9Sf
bMqccsjtzv19Eqooyyc9BlI5WhwiNdCTwXATCM1fpiKQp2OklZdMaGtOwDK3n2zf48VoDxiqm5Dw
XuddH2LiD+GZwAGywTto7SFF1wkLXJ+NvKfsJjZ2DzMZHw8BkoM3ZHbz+vrfMBjuUBVNpuURc15R
vKh/hbe1B2/I6gdiR/Cye1Qqqt062SLtfRkBLV04spxGuCknmxIv+bIhP+b2fsM6hrYerQxjssBN
9gxPevLXCtAkTk5ySQaFzmKZbUyko9D3zFl+e5gPkwMhvLNS5XnaUjy6ntoQPtevUqNLg3T9r1Lq
PA1jjhW7nf6Hue9rhlTlooOpeJRFGMkHQ2oHlhEzEQw6/z64T5ajSXdqutUjLNefWP8pn+AgUaLt
lHLSyHVFD1wDwAbdJp3+QnXBpKbCtDnXVDsNA22EKZRweFyvN7fTGzX6NqYWsE0T8LR8ZjDX/mxF
H4Hs3AEbD18mEka1lQIwE8pTsI1Ez/SMZ7qgX3L7JcOvCmj81suSZa42kNY7Y/ty+IcleNQNAZbX
dLgFCpK6+Q1Fgi7qVA8bKmKmboKNAJRrwxfTSh/Vxq5E4sGikfpKpR4qwU8eEmUOynB4ZkIKMywe
88dEKBnnDjRxtZCSV4trrmfCUZ1N4NRMZ1JqIadnDVJTR2ctcjYhNhJkQZMrM2p0niKoUxKmY5b+
YSqv0F12UW+aWBpPFJtaGpSNbw9F1vvVZv4wfMSsoQjr2kKQk78obtO2tVjOu2Chjk4qVnNOlFQg
uXFv44mqx98ZQfAw49wvJ0jl7E8+oITJmOPPz9ws/xG4+D5j0aZb8cMIFGrbUatTClve6VtrU6DU
kjJWWUdQhEjaDcxdpknTCNnkumAMgqReU+GpInKJfTRZIwhCLw4PdOcbjPy3+NInQMyCltVu+SFw
rMAlRKQi6GXTcQRaH/9nS2o5xX6o5UEH8ERao87f0b2LWSng/eF4K3mu6jqP+KattsWZhOSL3h8/
q3xzdWfkeuYBS6aD+RkaSZEL1hRYgnZ5qamQxZNQ44eomuF3NoDmAVmtSquGqDGTMkvWPrmDjrJ1
ECjFlYFYlkqX/bm3rs1kWyAF24jmARjlgmZSJe/dcjBE54LF1iwTZX1r6nPRnasxQliusvoXPYm+
ITskcOfxx80TnIBH1X74UMjSarYvNiC9nJN3HPyftRYmZF4TFcO1toUvIMuHFoxClgXzXySDLClL
4lWibWTLwXIeCZi6iNv6MZK3hhm0WHNJU9Sf5GQCYqSy9GTn5eaXw4Nrs6fZUv9UmtS81+wjoCKk
LmkYWCrINdvKUwZBrYCeVUQp7224T88F6DRBMANyPVZ7Fw2a6dvfMuUwA9QqseJJ9swv3Kb67aeb
WaPksywiAR1ryUranzDuqC1yUuL1EUeSxrJbBpufGbL3Ob1aep1pAxDgEBQkctPQ6n8E8mDLRalb
j+CUUwZ6vAA+kkZV+nvJLN7Q2u961XweWe3cgEh84iSS3KIiV4TvNZu63CQ+/ubsjcwKUUnz8+4p
Vz5EZs/x0QyEJDmsvrdh1UCBkK7dfOb0cN7TNdbHiRw3Tw+F+bsaAazYO9K2ppMEJoq41IOkoZol
gMtCVDb/ECH37osMyF9vhwfyLvzssB9vZoE61ETn/L3ZXQZlOL7tov6THW8Bl8hFLH/50U2a7KpC
O7GvjQgS1kCLY9ycJCvVshAs/DeBLF8zII4DWgQymQq2jfGHH8fSSLQKs7gq+TJvYXRPPr4xfE1u
fgAELZCcPSktyOB1Eg+jfzWFzBOSXnjjtSZf5aonyhMzuopAA8MiDoz7/04qdOdsYjv9YurFrmzs
BG0Ug1nN+32T7mfnjpEw2CJsKx6Kg15LxGSSPCKIMNVOH6Bk1Dz93rDSq07u0Px/LmGx/mE/yVz8
thVAkf8svJ4X/NxqwD5CJVoMBv2uoje0fXbMSC9a8eB/MxwMu3H+PVS17faYbC0APDKOt2RDUSPi
gCLbjs7yHvT7PmMCQ52LOb7BSR4ogbT4+OHuuyV7Ar7pYxEAppCOym/BjGrIfif1I/phuiK5ko8t
ocgsVXZw/3HZ+37hRe9dByawqjW2eS1gkCZVX357DrgqYC+KF1jwBiQ4dxizAHE/l17hJFGh8pTM
LZwlPqVtF8a+lmDGK22L9GHn/VQ0wnQwKRq9qYZHkqBl7vqd1X3OUTC0Onxl8G4zQh7mN6Z/xxVG
bKclHDdvtFEtSWrzssDvfdOJpis0kfLMYe+1cmv7/h/DORjao6//nBKFmM40q/2IwrzSgibBbUEr
4zJnE0cQtMDo74GkAzN2qZxtEx7SpawjGMYcBLrIz46XPeii6ON0S2J9b3+a2kvsF7dfKFvxPZZN
TTcB09JkkB6/XGWIZycVLeCEjKRxQaT/GAzQ0xt/XBYlT1POmw5UVyKBamjzO38DRupQfTsgYd4B
TKl93Jy0z/qfkHZUDr/VYCmQwlxy62kahaCBeixqRcCVLkQOpM/U69a5HKhDzz+9ULxKuGSvkK+e
Mb/QUVrf86axdH6zpJ3pAg2cajn0dol3E+MpVHT+GXdtnU33eO05fNMmbbhEKtlaraFtw2RG43nv
ZcVCeOqk1mg5RNogWM22XhhuhODg5jf0BI2r5/UOxUFqEkIoZNKfg/YmmtvThE4pp3QZmfUPt7EI
YosevWpqoJp3krAVX+rJIwd8Eb0+lQSGdDde2RP86Bhqunq0koln7PrhYAZ9gfWKHdIbes39oe95
MPP1PQJYNVFPTDOLvATnqMYzCIW8Bygi1elaZ1I/qrXPJ5C0R8Lusi2gjEp278n2OkHtWL9Q+eBr
/WjbvzM7lLmE03AKX7OFpD774Rn42MApDgmURPVJfK1gn3A72CL4t/XYjVjsD8GU7B0RPCvl1x7T
2gvpT1A0Kvh6rCqHW5CehlTNRVDgco7ejSUxXXiKawrY7DtFKm25iTgCkiC7gDeZxmmd2tcghWoh
uIFJuWBXBIsTd4uOc6APPTWKDF6JlUMPMk0P2UKgxdrKC+EOi5b/o8jaeLPjY6vYBYc9EUbM1eY1
fBIrG1UA6bkR2l2UYaZdr2hfONJTqVcXlVC14ojdXA/yw253vOYMSDb/QPAhxKCvGwHu6uGp6G/z
faV78Uq4qG5thitmxvFfrlJMiuYstT4lAC+M8/lbMBOeHj8xXWqVD2YSKErb03xw3hm81vAiWAsN
t8TlQBUtezXT6cNO36ba1+1OkKWdGPPk1pXFbIfC8EBnd+XaZ+xPdzFISnZ8TO6YhetmcdE1iFXu
OzZsMwnN1ewcsqhe9L3rp7SrrJPVsdenP8mFwenZCo0Y4wRXmDEtkjWED0LjMf+a9Pgq/qVxh1w3
a+wbsvTAulciLiV+UorjXDxvQaEsa/yhQPmoEhFC2GEOWAKv+saMEh7OQaI8zx0fYi86OzWqldH3
jVsqCAzN6/2ckO6ZRZvteGdpBXwH1hGm07jMieWdafzV0oaJ6MzeXH30TSzml0CdBSr0inskkVdS
Ez0NiHS5e6AhvMdOFXCmeJqeneyzzrd5fTEIiX6sDpbfkmeSnDzf3jZT5KQ9xiPlxuFBTpPi/cxz
5D4xoHisLy3wKpjS0pZEPkjBbCZ9UPHvOEbD9rMCjTrZRTH8KRdnCvV4h17wU+g0xooEsHmeXizj
gW9SVhvnYh7zluj5PdtG2MFN3aJH2fyX0E8JuoRyEEqUwnw1FX7dA9mFNJNB2NvEpBGLJAngshFv
Cd5jFsKX7P9sNeAPuG4TtJ4+/k22yMhtL6tD0ucOajTUui6BtYGQeTWKd745C5jTnuujjxa6176l
mh0nMH8k3Vju4I6ei++FkKL3ZLErQtGdeC4wtNCsV+dVRy742y+slxQ4buyWtdjFaMkZKnnztyZQ
Q5HdbmJcL62rJtB0qpXa3Crqgp+aut+z8Hh0eqgvQdDb5w6KWkFSweP2J8XU6JqecJBktk7HPYq+
kxelXuFfE/0TNdaqdRd6sktf59UgPpkwxyxu0VCCWoAR+XjBzVysgm5aVcoqwe43LIQKyC4xhpkM
Hy8pSmYBZqvRSRQCb6AeoMzuio5PwEl+7jNVN7NFsBwVHdKLc/M2xzoXaGkThdni1BgDVqr5hEQf
0GhyAlH/cAkaqxTBhbd3sXzuARy4GRJ1LelaFyYFLsYO5Xnas4WQOJ8dqRziFrJUVbvJX+y5jsXr
f2SnY+sIHXI8RrCsuepMb3WxUUi1aQhAv4VRGudxqONz4Wjy8ZoqmH8vFM5yDU+gjaUINFMneIRs
FKCiegkL1tFFJ/X91Ajnbcxd1e7pBl+Vsd8vAL/wSfLyx/pEGocPPw0o4DDmCKCMGryt2Hy0sIwo
G8ICCJHja5qbD2d4/cIfiA1VDN0i7+/7S3kxCCP1OdDahVDJeJHFt+b+wHVxuLbnEldvy5WybKLW
qifph/lQXYpPJo1SENMcg/X8bLKRSwVQI51mqlg+KtKHR8HfRzYtlgEsdKPbTcWt/rzXNobboYg3
37tQf1aLzV3RPCSPj/13ESZ2VF9fXx9/DjCKzfIVGFhQizexgEtAYoSEyj22IwqLMkAWM/7JZSkB
uUSHBPyFjhgIIdeIsstajcVxOux7TM4NDnjoQYiODnRpUhZHWBQdM4KNpyBnT9tWpQ0j6oqRF4Ni
f+0eCKQgUicUQpXpuUnsBeYGJG8dKMDQNvIQZ1XwBGxZH6jbL4/i7wF0E7oPXHrjTL/ZX2vqMIJu
6Ejdf9Ehpm9C/M7P4BeGrZ33egeie3gVsEAMALeEXax6G4I5F5PN8ioBNrUsbvhut+WfKlo5Pr/s
65RLcVw6Pn1AqENQYddKSGCIqj9C0as7GZUq+xCQajQMNKWaasllzWW4tzxltM9srZYEyXls5djT
dVl0+NvY6al8BpohygyLA4WJ4g5/ICE1Qckkp4alNc+dbmpwmh7Ed6yZlloRY01LlH+PmQNoXNex
GLQzzJztHq5B1B0ABkBwqtQNPubPIQc4MRTOc5K5mk4gV6Jd8a4lDrVEMS4T7O1hSpt/bpY6kfAB
Bff8gEYdBtPgCh7una8fiytzYQqQz6RV/E04bV/tNUWLbaLQfsBMHdoTOwOly5z3sheE3c6/p7AC
U/XPegiRQMG2TviWSmVnXhcV0GDOqFI9BbjivrtrsiaRxn/2IPZB81oPcMZfN3rkkpOl0MxybCZZ
HI0CFvZh/IULwAZ2wyXj8UoLRhcaDjzHZhZ7iQKSOYRDZe1EY6scmndpakznGMBSBXKGlL/myoKn
fBSpvVc+7qAc6qfvpkJPJ1Nlw/d5/Zia2Gdlx8D/WZQAKKnQK9jxFQY23wdRKcid2RjcGcbHkruQ
FrwzFBWpNu2CpfFUjFaznmj/caJb00KT91DCo0lvatNTXffV1E8279irdEuYk3WJL3y0peMTJhWs
yhG+pe7Bsl3xlBVCuPQbUUaivPGSHDPrwiJ4ZX83caIjajgaM+7sohrmv3nOuOJWG00kX9BlCXuT
/p9yXO3NE9jhwMN4QgR2LfRU/2bIqGlYB6++nXllFri5zvuEXgG4EtD1A1S07crHkA+2rqGW/jgW
0e+t/OoZBi1cfxitlNsSVgBGWU81c3M+P35OvK6jS2gUhn6KFVxbQ5tDaf0VkE7JlMkQWNtex8q6
t4M7G4KUuDuaSYc65Ya0GtW6aCRDuuvvRxulyKq4MSR+qtR86Yaaa5AB0ZcQXC8wQPwIhUBBnN4A
meaE8c2BUJufPq9WP8BgO/BvqPTxzntF2ZTRykWLmYtgzd2ZMpXzEX0zzfjjep1bNOzN+KBU+Dtf
J+wklPbz5HZKMV3rqYUb/szG3zMsqPh7eSL6bcgzte/T19/3jhKnVV34NXd1Bhmzot2NJwv+ZVpC
hC4M4x28Cq/MZy5Jd2UYmPx9xVye33ABpRUwwoPXMTAf+oD8gkx9Ujrec8MJJUkW/zyYsYzipZ76
hRbe0nKzwjS27EJgXfX9LPWcqoz8r2smWIrSMADIPN5iSU1K8QQuPPhwz/LmTIgBNIWDIkvvt+jY
70ShUCaP6VnoGB6UEORKcCfdHIJJ5UHlzzBuTAmuprxyLC/ICouTT/iqL/b10hd1UdaQoVJPAjLs
vOeop16ZVHkDa+cuS0qV7+qUQqEjv8h/1UtHL7VHnDk9u7VT+B0kxIxdXlmvS3jQ5pOxjoAvo+a2
6yUluG/+UJ8+41lQPFkITneuUZU4lI8t9vhQefnILVl9hGhfOe4O7oaoH3kiJ6ED5tiEIXhw7sSK
5OBM1tjcZNMhD2uUgp6IIbuvOSw376Ecst9Sa5+SlwPa81UoGfyXkKzEI1c65wpqPZ63qufVROVc
xqdKrUYpUDdIHM9rBPXe1WRhM4mOUwLkABw82xTpMqDXNOIGCXESE2UVt5CFsSiiiQNhRi03eShS
NeMd6lz1tbAegmXgOBOK6FFIoyT01otl/qGx17VTflLXgGVV2pH8OxCxTaHnLdHJzpzGUFDhi6VD
n9AnB0F1uJgdtih/TbBlxdWt28Tdrua70AjRKqahZKbG+CT+hPTTmECRpzDKriXilGxBhi1mEUWM
cQ7uobzvLf1+jM16Y6FgMsMQP8tLxHEq2DukfA0xRxofy2UIIScndK4X2sIhWfxh+bqTpbVjYnl3
/eGDTcSOCRpoiZJslX7sNPsli04keYtE4Hq5/Ga1ve4ukb3v+mXzT591sSE5Mc6NxHG0B/LE/jwx
KPci22ZEenMmdFxWZ7c5LLuf3HfTZzaGz6WiYh39WiTbYtaNxmVYOKe0pQUp8x4degg4MRdBVYa4
UB1p3iQYQyP+pzd9hwDwpNDx5dUcQPZuKeClR/7GjCI3WmiypNIfFBrY2pJhMXbm9hgLEnEVrj2t
8OfczV5fw8DLE+OSUgQhvKzutXv07QSmIphuisATZVKDZE4AhUTyWqQAVOl9/p8PTn4MwhaGMeFs
W8jIEMIRgIphkMWRjajgyp6o0frRkn0UTJyicQkCuR1E775quO9jJvmIngEMvUej6/Xgl8rj9x12
FRipc5ljt5p6EIK5Quk+byuz2urj88TR8Gl21RD2GsjKjnPH39qPT7iLABGFdp68xCpbwKL9VlQ+
QSSMP3ylrmxrEll2rIn0acuZRJTkgjAu5m4oN99lf9JN7/6r9zqDU8DyoLQkQza8miLlmEt3r7gu
0eBOr8ZmoBtMZA4NCNWtGSvSvvUB1KTL4N1vqF27wgsW/0l7rdAmzRXjBqW+n0vmaZ4zSsezkEqZ
GP1W9ZWl4UEnYLMhvsl3wP8XCS4cSJL/hcOHW/S4vE1WGw+d6oVstF/K8Z5oCwe4gmuSKj3a33K+
RiJ1GcOBbIEQhG0VJApAdIvnrcKxX0e3d2K5c+dThliRt6dz9wlCuHrNqpkT2XS3wUM9dUZHzbbp
L97uORjKiS355n6bnIOrzb0UuNUIj18XiuXNp2LLOtNTAJdQ9Y+qCUTdbWRueQ/0+dYS8f7KBvF/
yXM0Z8NzfPTB277hYsjr3N16XfI4KIbRqbFU3YFqDpFw7SdseWuHbKtpArJYWpZs1Y+PlCVeHePF
Zj0m+j3Elz+CW8aY4wz3UH0eyKe+Rfxj3OOz4QDwjg4w+ZM3kuLjx2yV6VZezrYVZg8iIx7U9qn4
LAkrTyODxHcoEa3StP+wd2JM8cUTCi10QgZiknkjlg4+3zJrHzLqQOs5vqTVOQaN0vIbAY2E6yLj
7JdRBzOaLQuMA+4jEEjNUmC/IdDpKw3QdjNzU7M0bXOXJ/jQ/z1y+d+aCbjcyaPWoOpXdkd5vFK7
E3PpS9npdeIVKcpleDkRqDvhjLUYHDOb1U3y38EmDl8IljQaj5yYe10DmM2ZBngqAadgjcqD+ugX
IWLjDwlWoGKqEW3S2+081MF060wRdSokTNA4dgu1CbTZj3QUv7tS/wTPp6/Q0o1S861qeWBAujMo
44O6a1W90/tf8JVO9oY3JS9Mxbb0gjfIqXnb0weDXgZgZ/PaXYAr4swXU1DokvfGipy00yCr8q4Q
5YGFexFsd+1UzjH6cVj7EUvTpWt90Flh+kbX9NEfphSHB6p7JV92BY04517DFISRhQmJ+TG0/lpZ
rrouB8Yz38VAtLLbSBaie4XYoL5RXhv43WjVFfotmzL8c3vuTfbHTWgqoRborOn0eCl44i7hgM9T
frIYg+XTgWcm26i6W8hf9HA1cC4KzfYUcYojc3pXXIV6anSDaJ+XmfbLFnhJus5SBxmCubVm4ZLv
ghGx1cf3aGOKfHaNrUTvP5OLzsezEy1hwBc+0AbSF8KU5L0zssxm3mw9AdTuGmc5gMoua1JbjtQy
cwXZjF9O1/1VryDWaRP+R7j03nCX1t6TdA8842EjlhBkj/F1F+NczfvQAuo4h/r/do2AipXzch5S
V7Izvs27ycOhB/ZX4rcZKBApUauH8k2mUx4qDRkm3cq64n+y5ekQ4XJ0mpIHJlaT/hOSrgGHZS/p
txaAXnAxQ9Ntw2KeSMwKoADs9XJsmZMC0nj2Tj7CDS2WAZEPkmwzEYJP3ZJ+yqN1sMQVXaAs1chf
9PqPd9myc5SVqwkHU0OfyigqlRnjY1pY/V09OLTiuNF4qwnfTDhjNfbhfAutVqw/ZbIjouLggLm3
9L/knpVBQuYFcD2t/r9C18/hXXsoSqAIVJGqRJPoSqxEfM34SApsOYVDv3zcFQR3i9HlJ9KTtG9g
FudG1Q4s37kowX+XPMVpIhUQC2JMyq7szBwYaMQZ3FeDr6ip+tONvoHOmeVYP9VzbbIe7xcWYZEB
8ij4UpTnUHtGDisZLsa//SRR2nw+CRz9qaOIgLkTBTkASa6u1rm/a4srJ+nA3vPK3xYIHhFDTWBx
dReNO57jIykqgdIzGcFRm1tffjQi2NNfjfJ7GLyeXOzM5OStmMzm1kEOIxkLgEuuvTkz0aZ+o4+d
QFzpv3WRzCPC9n7jSiwYNgs3IZ/bwF70AM8NhpRUczPblIkUqbRjmTSpZVHIAbYhzF+mPGP0nprZ
tgzktOI/8rk90QmxahOiqlnZX9wjP/QW7VxwxLPAIP3AeGxsx3FZb1Y13LkWxk4vzCBwQ+1NzxOu
tF9jzutpfGA5Z7djuQoKEicXL6IoQpyNmuLs6QACPVt7+2h/c+99/7p4zg9vq6zlBBRIbMj6MFFY
BEsa3HZqd3NLy6laotfcvdOZaApGYa4ImmqfIVdt30trZQl96GJukU9y5rKnDGJwPtKAORy1xmYr
dkJgeGFoiIHiQQB+HiF96oc/PQJ2g0KYRNVYbdwbOnDeUpeGNTeWaL7A8XoSH3amg6EEy9/CbETz
lEemGzDPpBK7OfT5TXDKbG1cUTIqO/xZ7yf++hB9WICfKUogx9AcDCq2kBAiL6TLzRGl7Xn//wTp
7dHa0KtSGTq96xnm9JFvX/fivM7OqrYg/7VYYnA/prk8RYqsVXZInXgfHjjeVDdG4/pYTqmt3IlU
Tbvf64QPwXJ0WZVehOhpCd/dqJNi8H96f6BIVLjLrtHd1jmuZxBdFcz1KIuXFp5ZA6YaxFIhsLaN
3swolZ60kp94MhYkmBCfTQyfQamKEqMAjNcQzXvL1Jv5eC3TnzmrLx17tkSS3AbQz8CITgPPn0TK
Rpw+ve12myYTogIJea1pz6RDEQPTb6inYR4GkfPZWsfCMBAjYpvpF5L5OhHOjjV4/PwjASCFsTGD
eBPiFxHIsInUDQaPcuj7pFucwZWt8ii3prU/L7kAhhxjRNxvX/S3SYtdWV2z8VH/rYwzczTysUrs
7IZQwvAbbR3D+JQ3GKsY0+y5JgwvGVQR1S7mefNUPqKDssuk+Zw0mV9c/3a72mCq6hiKJifGg24y
AnFoANsxZEZ2SoDEfXxp/y35z1ryW0rD5vN9Mb0SjwGeVU0LttVZvPR4vUU23Nq3pMGFtbhPVfb4
dKOucsJL0YxqLqIRzJ41fs1t8jRPRXm1FrcKIBR50FPslcSG0ef15yPagdiJlw891Jy3TnuT5tC8
Bm5FS9cC3tyvRVK7kS0I9lg9VDNltOoSTVF//ua8C95Ek9Dr9NwQPdlIQVPrcFbIn4FVVnqktX59
qSwq25kqYrSunEDgMV/LShV33nxM3iscCO2BD9CgNnRICZqpNSBxluqxmD3vUfgoPbIc2dtFRNMZ
JU9qqC1PZVsCZ0JSQ8XlACPkLYeiqBZ2Rg1dVWAemDmwcW2SQw4h6zL+C4wsn16IHwIBuiN2XL2y
uqyNDqC+iaTC6anuApc9yB3n8OU5CJNbPB5nGhA1kTGq1DA/KTZPql0XKmMCGUVeuLauOeT3X76g
+mSMpLiddN7tnbpiWnqYjZGcBz2HW34bS8o7a2IKugemUi6mBbqqlEgj3iZbNCil5j0PId8xC5rL
4R9bMZcRNwzfLtEjWXaMlkr+pZ3PWS2vNZQiJi7JB4SRrf0UHTK7eAedFib+FUESwBrkkktazNM+
tXNbcQMkSFewAJS2t4uotjoAQCoZ4XCAeq98fNTvp+uUrtQl5eZo1Z4Srhjfsh3LANVXh6yAYJx+
0NEWKcMGbCVI9RluBqjFoWnuWozQpDDGzVWKsQDnqK71Y3jc5tZYC8cD2dafjCCjUoqpCifHG2+n
RRg+iXM9eliD8eWn8sZqb8X+A+WfJfkE5jhNRfPXAJYTliW4Tfx1FTptPNURomhr3XbFHV5rkpyB
6dMTj0RTWVdIsprlF+IncUpq/EFw9hzjqy2JUFK/1yxjgeQZW6jm0hFpg1PIEVphdhLNfG/9wCJF
CqitnxxlsE4718WhuraBHNj4pdew7oIG/LUupnEnlUDFMWzVBZr0MEU3fURZ/253XZWFsW9Je/bL
LlB2/GFAmd/ULJywp7SPlNsiiUzkDkqrkEpC6OxUj0bHLytxU3+k/fIxsYYI+E4iZtDrRRFei9i5
mxbr8BjMnUC8QKp+FT8DFshjYPB0VwL4d9lMSNUcJUorfTGhvSvafJRzJ3rcBxZ88StbZLutPNgW
hlmYZWXbTZzVuW4ssa8xxRRJVDk+WB6X0Cz/2w7OFpW3+xvvNJ9k8he96XLjAjd6GWXc9pMPnJ5d
HYqQdlzWDpoXqm/9tTd6URTkp3qT75mCIqVCCT0GWskz9h2UhvdXqn8mS/9NqMf6lAK34P7uJcJg
K3VFFl2mMbX+XJkODkVUrM0AZuyKifY63AEIc/N4BtLIouMHmCIaamTYikm4LreOvU3+BuhjdoVe
ao5DYIdgduQToSOFyWcBd0dtciaWn7qhQMNUa9aICJmS0I4Q7wIkkO/xww17Bom1Db4JHjt818zg
fmTWZuQYIY6lAE30P3Vlmkrum6nFqBbWGnxpyk3Ij4LIi2ntSxsx9Wsq66k/EuXkNFGcDjaplPKq
hoGRZl78uGDRYa6vC4/nWPinzRdCZ/jviATrLSReffzBGtsX1qs0VmLTDg4tbNc+mPvm+LGzETIA
TgLmN0LgjHZRH09D68myqN7nITxt+ujZLaeaQGRopaOwEgC5tm4WgjoYMUmkpIpW9Bm68gfy99lU
gmxfvHW6jxwWv3b+I5ksG/KUFo2RyO1yjcAVE+IAzs+OJno9xmEafRFAGgrCJum77O4iYjhq0105
z0l917sX2HnSJBShfGiTUk4ZDIojldLTUlSLXjHvTTyPDKVJ0onT/5oFPydc8SlqLi4o2WcDPkDU
+3QzJYS7qT6EYrvOL3dFt1oUTND3R0vSGpxAZDj4hc29k9Sa+iz09BRUUA8XhMaG/5i6ihDQHza7
5lPQQpUjk19vl2bnIHGgeHJNWQHT9MfWcC0xgxx2oblkGJnNS7qob9xCaMOjGix8BagZCY9ryRLa
I+OvTkKcjmQKGj70OdOIJ2eiXplq75hdN37wAdn4Wqw08/+8LTsudD5BnxWACCCq0RBFxglVDOFI
yX7X08CSlFescc9DufrYzJQLlAXj2sQBc9fvPjD2BDstrAoFREZt/8yFVOEIHsmKhEVIBzN7wo5p
MU3/Yt+uQIll3d3H67wldFP2nPC/mOilpXoZqRyVdAiiykgB/NWkMlRYJx5DRBCsekNcz6rlVl3m
j6AUYIUDT1M7w4fes2RPUiZEG7+dPkp3GDL1e4EmJZoBzkMQanPZK6VZM3tBJ02Ts6fd0sNfR+6n
5deDi2L5x7kIZF4Llm/7aZHV/LyojqXgC8ybHIqL4GVmw7NTrVMYVlyQIQWtGBrQQmCClsDvPHO8
9MD7X/QHkCROrwK1c17LXCVx7f+7JbnU4kljrahVIFcgtUUFv8q41ioNdb7FBG6lImg87ByS2o9B
+v4afBTMWMNCDnxO0ogoQJ4J2zHVRV8y2rzOFjeZImnO44YvhQ9739e9jjxIyPhvj4kCR7APQP68
cEDVolZp1xwAw00ibeXBTImsYmtRuaBYHbWvbyTyZCXts4fC70B/cazXAsk8S0c/4XZRhdDPvCXZ
n8lM3Xoc420La7elcyqQqTnVH5NhgdpC6fEGINJDvGn9s/TrfadU/XQG49K2v335KyoxHLN6Iup8
IgTwIlvLUxwhxztrQFlhl7UH/OOkTSjRRypDFu3ILkfLEAI/TcImaWJcO5bEp35oRxtKSjpbGERa
kRqOR+ZRezmlrQ4I1/drw9+Kn0Tk/MHQsiYeKlW7j53sPj/6Z3q0m5Z4o+8BP5GCB0DEkvevMk6W
HdRk4KKFQzkStDh6wbyuOp3xkKXZhtBWc14rLEqtv9C+iA6WpfFxjXXnfgT4T+KfX1yrnDByI28Z
pwaGid4A41uGF1CaIVrT1KwGsIvMiRHuFW31CeIcJ9giLrHe4mYlcswqsPnksvKjxme6dmG9h0Q3
vkLvIJG1yd2dVVNX56HedyH06xd8xj0irim18qcPgXW8yupuY7drtEaBI+X4OkszXOzogqSAWZuz
tJmvk5VsDcpUE/TkA30bahzROcS5QaBNHlxcAF2lu02I7RzbVaaBJiwXdW3DLdXtodRBW00K9KRo
p8PQduGGDp52/WSd9e08l5LpL6sKZWjrELSZWpG7jkE6uAnJYiigU3MgauyWYCpw6L+iBYZQTbDK
ORMgtuExs65IuUPreCu1Vzl1KyhL28rfed+2yc8li2qn3pMjsMzCGRWFHwvUOg5VYM1aDL60Z4P0
dkMJ17KqqEDjTTAyavAhD7xdQ8O3ZdZsbYvWihM8MbMMPqMDr4P5Qjv9DAm/G5O+4FKz9AzqeDDm
5PP9tAUR3xCG9zBJbterbpaIdUyzZbU8gghaPaN0E/Yzrc+pr2VrcnPz9breiQ6CoCpDzQMNa59e
Z7+kpk1a1t7svvjwUmw/I+tHZ7gS+DPA9fROKjewQwJx0jdeglowmYOqV4+aCgQ6pHcML+d8SRL0
GzE3MpUdSJBUjOTCA4AJ4Nx0DqK/GYhgXCDwSwF8OhH6WX1UnUu7pYZrmv+5hM2/wlx383ti282A
HD5Ud2kxfjgp80KG2bHdqDrEpd235ETI6j4q+13OOd9Rguo1fa0MlY3mHY+WG5Bj6Z+S4L7AkfH5
cLAMPiK1l+0ebAWdGczTVHRL9pRF7z35IWeQ7VjjLpla87xGjjH7HA/0KQnYDdPHYJnnGA64KlBW
LlEjQCP1Xa2mtijdv5saHr6l8JhPSCcBDRJXuN+dR9jWhJwAcHObxikrX5+KzPuHnN34phHFxaT6
LfcDsglZIsgFSTI4jmdZvc9e4V8CZOoD/2OPOM4G54ckYqalD4SLeoFoMTylXVg2kr86PA7B3UgU
SB2tFES/4DpnKCORmP3vOY4aS/P5VU53oF3Xo10ACpGXu0FTE6AhmGuIbT+gPHKWgr0SPOkogqpL
U5QrtmZznQL0vKmNbzDJEqQR9qK/EUmETXKzy/SqobH6AXe5qL22dwL+XI0JJpeOnNYnm35+H9b/
iLJ7a6yXIouurJgKAIqznbubHUFED4QW/N3qozZWe00k/XV/seL6JWTJe0OlAaI/ed5dsX35cLSQ
o2jt/A2c1H3mLPBWD0xTPOIiRGr5FcoDqbiLVcHW3Hf3P8LehvDoP8ufcZI2xGCpD/drsh3ycqh4
CtjMlO6RGe1qdWGSqM2ViY/fuletFWS3HLtI5PUrUPfs3F1RspBT/gdEhe5phbFi5HtYk6rD04pu
z3jj1ncvY8iyW2UG3tI4zIOZfqG5nMoxBWU4R5I2WQs8t8S5+ykEU4Vp6BTHT7neZ/a1YUa+e9ac
gWi+X8BQ6wQCcSOG8oHoyNjJ4Z0hTl/DyN7qtEcr2thHHWXCtFAnVd65JIPqRIw6zU/v0RLYIm7S
1VCqMuI1fzHWi/KpVjMRPt+BRP0ifKenwoBFn2TDbC2GsnD8A/iTJ5E2OykmB2HJD5WLu6OIHnhG
gnXHtAsSRQdmwIyM9SBMAlWxPIWgF65Un2kcg9yxG8yaWgBN/zso841f/Xxpe339iPd0gSGQNQCu
lf0+eujzZKWFDJy1jo3lgoglP/uaiHYWd7e6WJDiH5R/NbJuzFPkKEmmzsCE84DKn5/JfodO8Vjs
uNBC/699Szbn70Y55hyy7UIGrcj1Uwwzdsq17vt7alghnCHAddkEDUeOtJ3GBzbqf3wNvj4/UOQv
bJAzMploZvXwvV+ynkOfaaMBKgdjoofN0IIVXC43qkrltXg/lomq0+WJ/4xz83iYrb2tb1ptNCoA
0hMNoaiiLEDRBmtWSuN1XcoUr4gpblPDnvzXRiYzABddSla2jvZA+GlBw1IoI3cHHrBOoGmY8FUV
I4Ma+10MnAOll37NOfmJZK20A8KND9GETG+GBNB3r/xrcMzS+rqcRVh5V3fitebpXUOUfMbAodwu
9iqz7CPxBgSGAAE64jSkMvbVEW041KbHJvaQ5MvJ2h4Rtn98id4LzQatrAKBtt2WTlgQfdJvyfSt
mFxAWT5lnBcAjXjqTIVPi1pALEmvNJJqiUxQXSLHtI8/e0mclYje5f6Ww8RCDBDjL/NLr1kGlAdG
KOkGWvFI//Hjq5X8av8ujCARJZBcAEVVpRUI/XghUPbLlRqFmyA7TewrJZ993cKblRpjQzJKSCED
BX3Lp9PiC8/wWeNMotKMRxhH2tEkHGzXJCZpzszAmid5VZ2y8QoQ3eJda4W2NbVrdygDLZDFy/2Y
lfuRDOb4rj4xgq11W/mTNCjeRvzCKdJyC8HgwKn2HFYEX45sVt68gUpOfRt7rk5sGKztXbXfUcGQ
u3k7KXqN/RRt8CRW/BV3cvL/5gBxWEqZsputZThGf3tnUTuRGIxLXCCRpkpg0gatf0L8/ncHsnqL
N9VfXs1fmu8ys3hEYfX88/QrzvetBT1DJpt744I9BDVZoI+kUamLuH5eSzjqFM06sPz/PGniOqVs
nLZ0ODoAhQetfFKDsGTrr8H61qaParxEoRgR9HXrmLSOB73Ts/Suw2qSAxGgd9hjQiDQyVw9wDxL
8Ie4lZgUELRleSOsXUeBC01kuSSMhzasm1fo2KrqbrHFxVhdxKZcMtJWX+tReiLQzJM+1QHs4gvz
3njwFEloFqHBy5NlTTmm+KvcTatfQDCTe0M70ywts8Z6z67RK4D69cGVvLk/OxgiVy5K5uAx65aY
ENXg+3Ghr0eMfuhN/h1izfwR5CxtUQGQ4vcKfCj6w2fIBgC6nC4jWbvrzGvdftwtl0vIIH43dnf4
A18sosJaFTBxU0fVPtlACkISao95XklHsq9QwFl64o//jeZtvGFBQyM/A3rlWe6CUqu5lpl5u7J+
/V5GXa6++FIWyhs600CmrcXaHiUhLzXIx3bySHMlCeZUonzV9rVjoR4gJqGWZ55i7z7PXaxKU9Ee
I50a6AVObtS2ZV4Bgd87uCLEHRlnyHo+ZcJl1lIc3jz7dtHNzwxrDfldnK6ZdNhV/dBdB3v+MOhm
0O2sGDt5xR9ten7iu7wtU+ZtR9ZBl9j5FsfvZisgJAVQ8/zAvkHxaLVGmLjzTRjK+pOMJHp0F0P/
BGrfp7S2lAZfgC/VRur6JwchOJIhAm6oMZ/CYlCyOVkRAHaco7QnSdupR0UCQ73wJ3DewGvH71pP
mesUGb2/5g9JAvxP46ojozXu+1L1c32Xtyto87A+BLrwtokWwuq+FWC5A2Wd6y+hfO3FAgBDazAo
1O00uPAdVhvNwLYdcn75qfqHq6h/m+dq2lIXG/TCoZ3BGqJ33SVe+dD6D3euMUUfCXtoldo7IsrJ
P49J1FJuwvg6QiY7sr3GKKQNqCdzzNadBVB+nMt8v2cT9PcX1UH93qKKlIgVesidtRzXnc7HpVm0
J2ZHnj6aTgXuGHIEhHPHRLQwjmljSFCDeXnpkNvqx7L3QIKAc5DrWSrWVyfYiqdoqU54SfNhDw46
E1X7zvjnG/1J1ntTC9/Lptcsix3MmWHYtM7KYw2GrPLkupUnz+RssBOCc5XEn5mFe6pfv9qRvCcO
pFVjhUcle79rh60bqx4ebrT827SPZWy5a7/whp2qBRhVMKbYl8YjH8V7yhJ4RD8fkMNIYIDljaNX
TEZ4dWP5Kqtyxq/eycMUN0S+hFm/3c+2kmp8v/+9EEJwc4y5j6QicukefQpbB2bnGwyVNwujvtpZ
Dnyv4kliHDOV5gQJ1SdGc+0Ps9cm0fFTuKfmn6PS3j5BvwWavtzDKvsfff4ELuZqWRyn2pCa8erB
yMJ4/gjqXnLb2VTAXbNESCDflRtnir1GKwayrsqYuPw82MzQS4hk+GeSqQQGQ78/ytEJmLy1e1zJ
Wz3MUJiuHlTGRTw3XVbAzpvJonWayuo+DsqWQtwjFNP9Qwv1hXkxP2zJii3f65KxzPtRzcTUPk9l
zjXgJq4NH95/kYik35xBBs29tH977ZIGrSaa+lwTyefuaFF1urcEszeqe/UIzyWXX9c2pbkeVHaa
Nux3thkHEp6c3h3SrXG8taKKEaYDGEMUuJ+Mmtu/V367Ct7GQsDOKOPYvky4zyqlXBWAa84oF+mY
cQ2wz/qR1RnPZGf8j8zjwa6iVmjJ5SRHjskBmgzOnpAR0ba/21lTwJf9/ESsiM5oHnS7KYFBxeXD
8n/tmz6oaEuzo5XO5SJsXji95w0OkJJcdrr+PQigmCOOQlK2+VUMnOeyzjzlaQ4e7iyftKNjuTQ1
W9gUWleak8LBJFHzpen+WYsh1oGU2xzy1J6eZDaxFqA9QorV4NsMKfVikpfaVJVAEIPJYLCbtYoE
OXgQJMtXTZ6/I7LqKAE6PMRv6ezxGtrqYnkFe0nFSAaUpj97IpLjWpCeoHqykiY7gNquHxo7tyRf
lEnYWE503asCWMQTzNLx2ZgxekY0vGG8PEd643fGl9u0IsesKKNuXTy5QLLwQ1JzjjqEfVBG0Ktf
BD5R+uqRhEV+qAlDxzu8UsaN2CCi6qvUis7kh18uNWcSD/4sXznLcr0nn4a+tAowAcCnzWnLeZ2p
UW7cH/kWDc6mXYx77JjQDJ/g5CWadtkU7dWH0bYc59Z+SGIhK2Z40Dp5rgHhLqS0XXvmcWmC7o17
1pZ8JY+iaPA/a1LP/WMBySUvNP2F/eIuXx6p0jFlUfYacWMOuok/WQY/Pue06kNez+Ghw8Mrxb06
PNv+xK4RBnYzu92w/0lGcBjcw9SLvCK9iArP1QF7D2HUEEja6f/zEY0gsyleLbRP7FcK44wICFSb
cZMXEQWS4ejlwWQJ7E+24S6D4qIquYiOJjEEn+8Ghzsc5wfjXQenRyjakflKePa4A5cWq2tW3guv
eLJFzIe7cM7fRm7BSMl04xd1krD1hkBeOCBvZcHNu4wOEMyoluQTRj43CyS9p/vGEM8twZkKLYkt
TsFlRORQsra3VlFxQ5TCFk00ljCy6MI14gqfbKBDg2H9pBSF2El2GAxd4GAdJS7zyke92z0MUK0R
NlD+dikLVroAbXyZAlAbVyc83AILVIfcd0NSDp9o7HJt+cUyRWDDY1ARAf9leWyQTEYda64bEReW
e1lZCZOmmdHtlcHzL+CHVavYK1F4WuyWjJfrysUjzDjHvVXs4+KHyBRUbQgkCHHO1qDKR7IqdP68
xFqiqEoAN/BNcdIRa/qfd/Ph9jE4a9HCSIoikKI+R6AjM63bRLDggj2w7IMlR2gIPCXDb8Ush9mO
zHFf4Of79ZX3fFSxZ+A4xprtcI09JSECe6Rufe65c9M+IGsCEpeeqlrVylfkSYFlS9ZdOmxF9BE0
ZBFt2PKvnFlmtY6h/UTpwmLQrlrehk0C/SErA2uzjkrFvn8aa1UG3J6U3DqHZVzMHvJ3HxQ8KkYr
2f0hpgg5mvdu+sjYrPbPC21auo02hM26WHaONxwUhk7Fad48V6nCNs2gvCyQKyxGd1txhcvJNmkt
PRDOrxiuYq8L5R2sM9spVoqq/mhJoUDGstXISuHEZHb9muBQAxn7lhghfIU2+WOrWmh5Uubl9CIy
S4WzlE3RffT7ScWXRqgkSRy346x3s6iN7RHYEW0MV1+MTTrxALHYBLeL8OJzSLf5AXlw60p9Q419
LlnuuYwsR/1kvch44Cu3AjefhrwMZELDgDQMnlHqwRkuYPzQB4SXU3eix+2Z1Qg6Se+bDpRK4QHL
rmfHXv+lUHzuAT7O7aYqF+QVzj/zow3E5+T0j1IpL7FdOgzU3QJsv6/1N+tnMIoKcDy7MyhSABn1
oOAUnHntuda1NQi5A3KmbnSyy6T015TQH3AdeNm0KG3TQ0H8UYJjIMqGSHqgift37U4TS6vpBQuw
Gth9EGxvECmiZG+cqGcAWGpeUNjVfcO9iVjJb3ynG4g2lKcStoxi08P+7pH8l3nCX+7frBKX7SrJ
lklhyzOnvjvqODV3UicWCy3iVzaB+RpY+4NIVdCECoSeR3RdDzIBy5Ft2bgXbkN5/REu2vHVI/h6
KQPRZVOMnw4tQ1bg9svW+vgUDkpBPRNoDnsUIMgyiMlbwU4HRyCDBD6yC+ebaRW/xzKjHvjtuR9l
bswMwkLqGNEH/qFYn1o9RMbgdGNHjuFDSSZC7GJgDAKvDwxv9QR4yqz+UE+7IAEFc69S7shTx62w
19dWNuLlRv8dFKIrM0OUs5RK/RxzRr9v7IbYYVRNuTgaQUyIHC03VJtaX2LCFHzDR6KTB+pOK+BU
kkl/jHQhld3BuimyYwOFL1K39AwkdG+ARlKgjNfnBEqzE0V+dm4E7LawJgjr86oI1nyBvWFcgI5W
/iMmKR47mEwX3bBdqA0dQz+fo473K7JuDmV0JmBGl5v4eOg1zMXkB8a2iHcmJOt45+VDWo9wxP/V
GGlfR6dzZeFI0PgvQWukSa80jk0GQjyB+MKdADR+unCSgRepR0F5ODq4gp26zKShOhYjsMGbxC+Q
FNdhNf2OkNMliUPsJ/yXjzf2/C7GxKDHniQrqdwpryxpSkril6PljQ1DbMwCDofxgevu+U3W/84W
nvbUzw/mSD/ki7p3F15uARu3dHSlpIjQoTVZprRX3fP+I+MF5EfNaJb41vkEBzgy6MIPVzqWckQM
mopSZZUB5XhZ8QnHDsYmPUX+f1NTzo8vJn1CfJbg2syXI6QrrD6QoALmOWXb/ddsrXu/K9En8g6T
voNiHpfx3CzyAyVZldelnb6iCakiOXgYuEzxtZ7SaBuaKRx3uBvzdgwXcHlvS2fUn+fd2/HxF9Ee
jIGx8Awnekb5H6Tw1ezjiXcexM+FL0hNPYLvxIZ5J1xl4d3E4rAE/EkyW9sBQywrlWtDWy0l0B7E
RiDKt6FgErrOnRWcc9p5ynYuxJdobdk4VDbcjY0ADqkSAu1j6hV/pdVLRB8rblMr4QphP6Z/is5s
enI+/ntjr5D71Peq3YsQ/rZsuUx11j7KqoUx4FmIk3JdiBqG6xPyCq6WGGmbfYFXyKj/uEtMAq2Q
Ld4tW4l5kqzvh3Ji3LBW+ey0ukoxnj0K+dZktC+neiAMu4H7C06N+SNXw9bq0eBCxrIeN0+8ZUII
Aj2FVxCdVunFM0onzdNaHWcbkSP9TgoZi3PMrxMzMN8LOMLbiik1HDavzHQgb/vwbqnf9qKVT5/R
olgApIRH6GnHYYDd+XDhYLzmga2gLp3TGk7Zs1j4vj1t5jZlqsLXuN/tk60Ce0gqb+RTp2yn0/xk
0rEX6RCbeb60rHD24gUvPbFM5z/DcRSbe1LY8A5+NeC0dwZeYchYtLD3H9pqxVaO9DclcHRLniga
K1+zeqYbhbBZw8W80s9aM8SMw2fYR9KdXiqU5dXYeYmH1GfGZXgLyqe3V2i+D8BySJ1DTMZYJtxS
GQ8tRGInC8MgsQmcruxIkhD1YnaHFfGG5x+1067Il0Kw9zy6F9sTDycAvCI6lIkZu0mmowXOp3Nz
05fQqt5tClshkWDt+okp19J5A45q/bPgCBb4hRQ4GoqoNypHsmgoIUoCfz2xxB8oUguP5wvik2w6
EonKBejACZ+uZt/q3nD4ICYSCmR+XAQ+CiFLKhK0JuZtkVKxJ47N+7tCH/dsh8JzrMCRKxymN5VY
1fn2Q9QEG1qXjTbfCa7A23oKVRhK/jdes4hHf6BhMKzMO3d74kRh1MJ5afJFDNsfjveZ+hWhLFzf
MAMOBZE8WQr5/3SU0LyroipNF111wwPQS2+BOncpeQOW7AEMGYtkf2PMJ/RXsBjtG6soM12nBt/x
xBMCthOEw5cywXoo2LM2ZzBuYHrmqk6/KhwTiS6WayF9STKjPBRNpRLASirCtQ7+PAjCStU9zgam
9ydjZldm6wO+UqDALIApn9IJfu2W3XfvKCtpQ7Dn5yvp3pHA87trcQb+NwifhXzh8h5tf4AyScRo
PnSbF4rH6OZMnOZvaTHEc/OlSli3yFBpIwHWGyv216NKWJdXRjZ357N2OR1ORgrlct/goT890e5q
gk8bP+yj7HC9i2uNG4re6zCgwJOnRxWfnGErhGLNsNr1kGvKusdmAiTDivcoB0a3N6ZvE3WR6b/P
MbthuMvX/auWYStHREPQ1bt0a01D/kHYqaE55PL92zaFHcZ0O3gb34Uux9JD4XHaK3kZaS8lP3eR
Jp2N+xFQhNvH5Ti+AgSjTCCHXioMnk5BPsHR/1kpZwhK6aaFGOrP+VjXZ3JEZcdc4ivlLjkl8KLQ
h02B+pa1idrrvNj3LmvtBAvgHno9gBGoQm3w2GAb7Vera6aNH28o+4o5WtrhGE+h+7kqpr4Zf/lt
mGQCtPDTBpM9377qGBtvW/gRWsn1t9BC+LXUiCXPvAUxwve4roN5DdM6L/5uTpw2jqdulKpkP7GB
V2uh8+tXmnM5c5AbeD3DLH8X2GO6gYNwJs/MDMAoSI+YMHqlOoh/f8iA3In1HNsMCM0AH+GxSqie
lltDvito/9w/XSaEqOU7S28FU1A4vE3pdgu0URw8fG2H7yzBrIEqLiBqco2NmwICu1BSiSd7u9JN
nXvNBUbdbH4vD04H0BY2d+4pkAvaEFCJ8kyjeNbk+9y+r2CX9Q4jb3msD5UJiAFSnpoEGfS8P4oC
Vfcs8VnkyevgG1aKy075aBgTY8qvZHSZkXAuYj50AXcOmueG8vU/MIlx+OzB0CLRWliQPfzfFYL2
o6KX98alPxfqwyEyKkjV0TYqSqegkwI579Hijy3nA9AcpgVkkwcXw5z94s0pC76LJ+B7A+9DP50f
uJV+855KtF4F0SLZxiB3+VoYGf1XOxq+GjCTX459QdT9ok6diQTEFaM5kc1crSPBtaH55deOmS6A
zdVwCgbcmJGixfTgKYncYpsVNwNGxs3iA9or4ksH9oLcKKejpt+WsvGhV+ucnZnGJg/f6WBeeXrP
W/5E8hNGAcwNRln5/ThES6dEhhn5CB38NxMnaqSd8MYGE6V/vRXVA9xuFsf6Zz47oM9qHAupb7Dd
KWS3jEhHxWyDDAZ44mmkqqZH5l1ak/QXiEXqeS9vn1Kf2cim051b4ocm3yU98K/QLt0RjntuOrys
oqczrnDbRlgR/NF1vwXw2S0Qo/lcfH/DECWxd/52u73Xd5u4eiqPYPZQdjI6SIWWVstouLUzkrGI
z8jaWBBW6FoJm7hOYjMBjY+NXnMANgnsRmRmAuUrScmp/isBxA81F4O3+5BJvwsRgpgSRC2A3Ju6
McgisDTttM9bDUvCs+YOHyIHUSWnk3qp13iZqRKBZCZrGBBHehdtcFheKMWDuiAGdZXVVUNL/6Zu
/IC5ZNe+qah72oxiyWEHHq2UYISnn6tDjDzavFYbjmZljvlTo6fyDOv8mobpqMsXyi6y8EUozVGJ
IcE/UXhdBqyywY8Rmz3voeMXu1iirI6rzfYS9t1dDyWC11kefDSHQPjE29/dOaEz42z9rCP1766w
ZnDFJJjfBsHaqSPwT72CRxCjpLqHQ1pszdpBY66a/iDiS7ceMteBpCJWsG4yebqFd2wtlJqo7vMN
xnQFFXTZOrLmOv38dzqToBftRrdGn3DOJgsO6C6qQkm8DberZ8D8SAzbEqePCeZqwTmEzpK8pTXr
c6FnsurkPLbQ+tHNfLP7U9Dmvdzx6k3XYZiFOw7yfdjYOJv428mcuL7UvZmcWW3xkg8kot3mgeWj
84tf09LrC98C47199RZX0sNnXgeL7+gKqnWlr7rBWHTZk7mYgDcny9Qxv/Z2y+Y29/DSM3f5AVLD
xOLIaF7q62yCkFHJXqPemDggncSGwn/HTpNiR0ZT9PUHgGqbseDegOjZnFb+6B+6lW8Ps7KATA8J
M7mlLJn+9Xq9E+4F3K2FCi3zTCr7VrD6nev/BSomfuQLhXsKP3HY3zAOUPR8UH0Ds4VVuE5Cvrcc
ebVwXHxaY8AG2POVYtG2EmVESP2hTO3r7geQ8xa6Pb9cSM9VMydadOtkz+Snj4ipHi0nuJv8a2I3
AAlTrr7cJACkLHowV7CWX8aUU6Y6esh5KmnHu52V7tfoUBgsQj3+COrs4NxqKEr5lLE9Vq8MHHAR
afIvqel96sTL17oTxybFvNospAqc8xMqQ/Znvgse8h1287HjeKI7fIJniZdRWbUojZtdFovCk2Yt
C5xgWDd/0i2bIowk7QkHAUymJEJKc+cpI+PnkCKT/nIy42AXWxezg1MoRK8Q7Ztrbm/FHd0oSkfU
Jl0Ntcoy8YMbCQCqevFpVfI4xqUMGAs4CLmrGZlYjxSfPmDwR1pamsyPf2yuONg/IrsZn1Qa37kJ
l+j6VaPqeUpyJpfuK/SpHNwnIg4ZZZen635NB7X6zY2BN61yxQogHgcYfirnDT63CCk/5XioP0s/
GFgdtTw3BPH9V7ppnZsSAukRdAKnofGMwToSp4Q87N0dQz/31CuoWBn8FBpeL1LPmm6Nqf8qP90u
Xg/bUkC46ZPHgYqSx8V6CI++KRUG78Z0YSHZ7pUFq+lteduKoPiCXvdWPV902bhrXIF6ET49zO9A
Cba+aRZvW/V4A/SSIZ2GcpCCkCJZAKKfAoFUzfnBTkSEc/44cM/dw56Xx63n1QhHoWIgVPqvDyDU
dJOruvU+JzUJVM4ZDH9N7ArSkmPTdj8DDCQo0nWzMrDeqMh/igBq0m/k7to1AGan7Tf/AmLrRgm2
mAmA2a9mCoIvTSyGgP5fpTUdJzU/iwpqjtzrGB93h75ERWNYOqQoNOrtDDm0tXvRBim82fZSCw/K
zvFxc/0ABvpvQ0E7/0E5tY7oI+gec5xhUx8kEkEc//qwoBLTLkQkNXko4rNv/W7NSa40Ro9WZmmV
qJDeV3i7hMUoFtt+KcoVisTA5ultLWPr5Qeiv2TKrdkQExe9rkZsyS6wwA3/hK9RVv2JaVaERC2x
kLAFNRZly1yhyZ96dQ1+v8+SyuOGpy87vEkacKLWKQmNsXmHLPq9n94iDGXJaoFpXO8O2osojJlJ
o3FtXCnyB/0MlW6jleJoz6XImAUIR+EfYue+jQ8D6vad7uL5J88UYlSlKOkTlGSR5156PiQQXNbY
6zOOk1JbbxQB92t+mfagK1Ka7w2nJoiKF0pPvIbSx7XfnA0PyPcHdVjxYjzAhE5kXiT/Xe5duwEd
EIGHr1zjHCUXcj+PNLh1zIzKW9h6o6R7uIMnnaOmzpVox47TzzLQQJuu9uQFn9uwxFayEoZLHp0a
SLspwczFAbmjRWv0qOzn3mmptF+Vuw/RNpORQhiNAcOnOm6UY+G6ZJCNxlRBEECmD0QYbRAkwl0j
gzXNencm7y28zc4myj6jBCe+OnCyyVriT5eXqLhrUqqYNnCkCdvIIZ751x93V8aAGiyiYa7vvQtm
phORDL6hgydYPT5AmPqw8D9t/wzDXBj/aGvZTkpXolwTgD+8TsDV+slFFl3eUJEKybJmOOqoZNh/
PSY++tKdFy28h7hR5ulS2Djlm9X5hxq2XH0zjRmdGyshhyr4Kio/RknRD+q3ZmHvWBM98e+cK9fa
RPnTdeW5q4W3RhW3lH0c2k3Hhe5vjRpKCHFy08JvGC8fYMr0jpZK6UCVqBWwfUq+5hM5ywDxhGNJ
86yhbi7RaDURnoD5M0wuDf19mLlfwnXg04ATW6PPZ0ZsTG+acy0y3BwyS4Dj8cLBPWnCEIWaCX1F
bLwHP3M/AgTtNajqbLgfAMpjPSQzdhcPryfu2u7tiP7aHfcimsDeJXFNNXW54L02s6QPKgbRzONQ
1PrIVSzBKy262jNrRTv+/i2WSYqc/5j4UJL7OTwbgM/9gvFqFUUBWRemXdCfD1irbUnVVJxBq3Uh
Pozxl8EQnEtX6vzdtIHQI+RRzP7H3kbA83VZYSL0ACHKb3tGsxC6zWgTsHRChUXev7MZuQlt3y0Q
R9XWPR0cT7BAAKrMMBR7Nq7QNVx86nFwmDj2D1T8CcuRXbJJS7aDuIv3pJqSEsGT2MxeRmUYZK7Q
6NLFKJfV0Nt4Bf/BWc3XlzdqO6SMCYM84gOq9WxJ6Z7qSnIVXgr8z4E2Ee7PBq+b6jsfmqy7hMRa
Gtt9dxbmcwVafuUNRO6IwNhEszfw5A334mtUPm9BINjSTE2Xn+kM0BAMwF/0KUv6XKMRX7lHfq39
t2R4SBrwH3w/XL+4cMFx7NObW8YzsKrSlbrm4JOn7jc5OHAopeMDbcEz7j4nEd4eWGxCSrM2skIJ
8eK6i5kJGCBivLRXQ9eSUh+C4xmNPvwNic9/j8cCUSEeMZtef/5jcf4pBwD46xbiNJW+L5PxmsCc
uLlLqtZDqNvc0yrPloH+Pogg5a+Jc+20g0c+z+r+S448xKQfcQYSVOR2edSKIzVtqE2t3Ss80AK0
qwT42Ll+xIq7Frvwl45nZqehoXtiH8xlzBSPB3Flpzot/Jy1+vzFvYiz4MZC/FJVFYECNO3cOekX
fVc+TRSODoLUtLO72gUHh9at7ZIJ6SfLsT8uYGrTeDejYTy/XBs9FU9VoGyh2EdF1dxG+MkyiS+M
tWUiKn9OtzR8grPctmbIrsoHbf381rxXvkeso0fvztS/PM4+23lVuJZKWbni1PPjAH26UHvGeNGw
dDZWqaNGvSzqCwgUmQDm2wh3bg2tpdoxww9wJuYisze2jUK6AX+OEoaCB5cswU6A5E04i26yVH93
D8M7HSrYa+oMZt7NGgb59cAAyPDXNlGa9rQklWFrzieXzHQy9PrbQux1vxEaVYJc8w5RjGqkAJ2/
y3s6KmmbKNghx4e+HNszO0RwAu7rLlTPF9cIemgoYxb5ZRbuzM0apx/E01RqnNoEJH8FoZyI+j7v
PGJaQcwaUN0Eb5vt9pBIrRn7JuWliwUaZMAVVLUrVCHGl1WgBs/JL6fpsSXV9U89rs8yq2TwV26j
j+oR0MrjGdvHKr3wCMplx3Zj+wFDNhnaV/Xn5tIUPRKY3UdsBOj3je1jUXIOg3FzRM9n15SRcbZp
FNDQ/jAHJnrOeR9BmEOImgvJ33WTWFG1TRs8dNQDpkRfknVEC7PfkXiHDjtMbDaaVA9nMtRBOLrv
dVspOeK5I7zewqJsjvgnGtpADL1M9lXqAow9gPp4i4js+jch1b6WOvEmJ3EXmeKjgU6QvitooGRE
7w0Hcyt5X2PODYS1RT2TOiMvTPlbuFlHiBxa0Km0RfG3Th2EszQt6ZnWUj8qbAtVnsEfL3O5GjPH
9y5qRTQXiQkeSP1GiO2kYwpfRYkchaqoGHn4AxOb2jLy7KLEBkevvle0SEWZmpUJVB3Adpd3/1LN
yVOkHzbH2ZpsW9WZe87wBm3Jnbss0Nw4XXhWwFF1+VDllqzsBYhYdqeDGYtBPyuifbw5selJITht
lNf5lxI8AvMOFN5bFkChi67HrjMdxpZTfVs5MsFUn3S35lqkvdPafBl0AS24pwiSUxF7x5cM9xIA
IlvCWUKsHEC7Y0bnsEDUci2W+zzlKb8QIibpqkgjS5WbvbL4VD+MoCQVfyuxThake2iOqF6EOPJf
uIEo51kLuvyDgjFsB2/EbAIGBRPKZEWBuQgYc7TQ8YusbWQZ5LxU3btojhwosFW5GLUJdmseN2yo
d6EbeSgCw2+7GwIDJwM94ZORdE1IEwLEq7R7186Uf5dROXhriGprMlSsVX86JfkORGXGCjWdBajZ
mw1QDOpvBSMzfo5Y3+6c/8Cs/YIrawDRugKAss2/uhkyKljIip7lO7ro8sB+rLVWsYEIZ4m8Nl1/
fwRAcS8+2UE7EoMNhkJz5D6C1HXvNRwc8rw9gGnjx3SdzRdkv1Z2EJxD4HSp+yC/zHKwJoastiqn
VUN6w3L7BbBs7xXq2MR+ceMuNUeOkBgrO92Ik106xB3mxXvPo49uAtVilE9uegFcDfFMsr9cWR+j
0DpklHA0IUcN/ynXUgx1ogCAGhEDl/Pw62JKzOnNIOoVV5sRS7WvN8yY7Y6aa6rkspXvUe0yCApP
rIENose2h52xgwz2uudOd2a8+np228V5ehvfFEcAdhtzjVFMERWzQlL+mw2LeC/7B5l9Id4ick3d
e1sNT1eDnsc7XtVxvOZISFRinQ6423S/zZiiNINdQpEJMxl7JeFRXXIV8blyClaD3raNmRhPPW+T
aEwoyCkIEK+TlM8sBlapkZDiCDvMgOlsJo5vvBPvglExL+P9qIZxLtrEYGROHOKQr2Fa5Z/Ic4fK
eV6or8g1n5uYbzmMGOOFIclOvIUBr0+5+aYZ/NzmohYnOonjimElx1xRjvzurClEuAXjivM/BN2w
APTm3bHFFBF6WG6/AG8cRSFnFYRua/3RAjDqOhBRyYgxeYb4liekRw7pqa4XqI7XEYZIsOucQxNA
tpzJBAwpNxedwZmfcgi7Y9zG8BSCbExcLEn90+yJs6LFMVlpbM9xKRZ+ZnF2Bw9UqSRMKgIHiAV1
krQqMUjOLGTA3cW9beEnJS2p9ze+418O9m5dp6r6qNqwtPYMFnrBbe89hTDdg2MF2xtOyu2qAq0w
06BCO+5aOshJI3ySD5lDHt2MRy9iHcA93Hqqy6JsZvRUG3TbOEw8Zu5JuuIhjVNkV4B/7AakcQkJ
kOYFAloGWWF2fwI8y+NFVMLoqMAV68me2lhIW7kcG89pibqAta/QlgG3petQoApOnQmGVyXhSUTS
H3W0pQziSKv+TKjg8uH0vatPktghKvm7P7Nyfh9rz0LS0+KSTOWsU1i7wx46wOuD0ZOFQ2Nj9N0W
bxhZuvpXuChJqn8rcMw+mWyhkkPe+kbYdMMipnGiFbmH5NS1gdCHzowOtUamTRcN9kR6T9u7038L
Bu/mGzOpnB8N+CgiEFxs7rvDkls3Nm9a7GTQkimOhnu7vEuDAg+QdUAf/l/8FsAiG0U7kLQuknW5
xYjT34bOzoY7viLCB2qBOgUCKVvTP7qTa4M6HcDjjqdISd8gOsVQnFIunzzwie7VzRjSwfPwsA7M
C/eA0jFOw36En+TLV/zB+2pxaXFfHtYfUjybEHf862T3V48VnrJtlnuuzMfPyb3UxtURs/aItyIS
zQ/ssG7oOTsjNzgQFZd31MVkxEmDBs1lVN4oXwLxdVbbt8khFV+nWtwuTQGJRmNpnkSM0M+Locgr
PYy8W30z301lZnk1vbOZB8/vP815HXRr4ybMrkmeVJJKot72rqM8D+UABmAvwuaQ4vbAeAOC1ocN
zdZ4mbYp81df4XRmaoQafbxuYOqGRqZjKjVc+yQ1SLO38i6af+C1JPhQcx/SX81MHxXnfRGiC6gc
4lNvVZH43O+A+a7/nnk42aEDzRfVFi7VqblF6K4wA7/3qhoB1UJhI1snLn45ocTY5wOWelzxNhv7
IxqrHsDCQ1qoRPX4WlLtge8Jg31i9HXZMv7T485Zdgj7/omXebr476WAlJr/81g5bKEVKI/lpUge
KWNhdD04IY2Z6NNZgYLFjuVae0zKlO+n8HM4egA9vS43HqBSilatrXVzMz7kJDKAjLhWbO15kmTA
y2LhxIq1YFj7JX3DISyXKjG36umnD+/0oYVSif6AmQTd9eCBf7LtNT980APX3mgJLWZ/KwTt7sAy
8RPYXW0bJFv1V3loloY1eSdipU62l/Uc3SnOfT29KUqxG6FkCXryQ4kjymUD76NKAkkaT/zqGotp
TecW4eTG9xdayPyu4eYcSUpOfeg2fBkqxt8jUAPzKpGFLReRxqRpZRwwh/0qW12z7Z8I1SiVW70L
FFcbavvhYlqyzuPjrOeAIQt1QZSvbyweOj5ca3x3Gtte3vwfS7KKSRIjAEvV246zXCsQ/Kr2x+Q9
Jw+oyYVJtn5NOiPt1Ak7gcC1q+P1z4KftFv4HRXNJGjycq8VyhAVvx0MS4Sdv+qLeBx7e5Uj4jIM
gErs2ejkso1o9eR/X8/Db2Uj80BMMST6dTRPYWQcwm+kv/aEnc1HdGYnjTYs0R7cONRkMAH3ZzMR
cyrkPSgb59iSdLtLUfscuSEj9JmqgG5Qeuark3Mq9rsENxYthDSPeMqx2tvwK4XenoR0hgyPH5H1
tYGw8xg05EgI6+IUuMeIgwZAQ54s7LT55P6WUXChHvxkxrILOwcoxpT9vqHJYrSpjpR+dqgOtp0g
gswdNERsXTDDqVl3OEyZhlwLA+xLaJLGWcjSLlGFjhwJO0So1kyjzW3gr4LOr6XKDXQI6WwnAvLd
xRpFOLrafBJSWS37G90t2+UdmjdMv5PSjzUTc+GoqAW4weDbaw5AUnEgElG2/Jgc5waXws0v8+Le
XcIm68qK3qfWqnVzxxnj66ccyXLgHRnOt4eDbfSv03KJfn+52rpqRSW1noBQcuUYmfNm3mCd6Rgd
L2VANN4EFOK48WA3qDNdn0kzrxN9aupI/SuQxsmlWRdpfD+gV1CattmUCbTlLbsbeq/YYmHakE0z
LzVHv2XHwwVSpNIV44jFL7VLsh0624vJ/EoTHqUW0A8HRFKm4rUmm6FqpUsJPVedUpJdpnj25UVI
q719pMfsDLLCaZe8Ohg47KmlF8UHzplZ84XKyk1JcS4u9a/i4kF2bVLV0WEXS+EIzZbMnUnxlNe2
9D7NIUDl4WGsnc3Q52ydTaNWw5qIb+0vhqoQGdFWM80Oukc9TnOdy7Zo6l5dH7RfyMlOj6bPCIO/
VFQOwbW+sMHyNGuzbRuMVUI/9ytO7aLGk5kveQ0IDkd+Sr4Da7ZQY0/LCI1SE+KD0Aw6Z+1bCmxp
9UBRcb0Gl1455VQ4E9AXFqTLBb9qYLx3Hpi6spHY/Y7br19CaZAaZv8BXJHWBunX/UCwhtzhmYUj
F3PuWboeslk+Licv9eaCd8PINeS6L66mtdRIt0hleRKWwGZI/tY6r41EusE8laD6Qdb7xc+0EXmv
7QxQnfRn4WpcsN9E1pUpM2l0Cs/19JeuE+/V0YtbI+KR2FbHAD0fS4TC6YEPkeT61aXYYu2ktGYU
A6D70I7XBRDU+KS0PX1CmInY7B/LzoIatxYtcQHv/rGoyMqhLExhxf0FrUbRzPwgny790a0zLwul
HsicNAx2TGJG5XRzc7rum9WzWFjUi4Z1wCw5sP7+uCNPG4KSwCkPpskqFSabP3m4Fnl7hnsFtL42
NS5NJ0FQyxhVs+c7so8vqBx4xbhLMCJE7LRWh5crtv6QnR3dJ/wHTQiDoNJpWThLV4F0FFPTeBSB
Z3pxcIjI3bUtGD9NVC97oVHNhTAQC1hxhXQuZZJ9csIsYJPgjCAE7QtzkcQ5WsKr75mP67uEu2cS
3R/Q6sqFEXzfCOhC9D8tksLCieN52a7Hc41VaIbDPW9FlPzkWesaLPW8ABR2Cea2pZPfh2awHa/Z
t7gWoop80eLEudkR6TVeAQdSWrmAlA6FS43UB6Wy+GP+VgmYd3itKjvnPGzAOJpiCED0RGYKyolz
0CrDvAzBDtXF7mynrXZeXb1P/Ot5sof8qt+zll+VPdwLEa6Bf+Zuks4Rt7p5jT68ZYCw3lMxtNqP
IYrNco/3u4GuD9/vc0FcDn0yl9JjLpWptge1nnKxuJ+lLRFVcjeg2i3aKo28OM4eRZbmYsN88COY
y4DiokzR7lFHLgEXaBDZ4bnVw/obxvvQSypb/dCVdGJZMGuf+Grmp7GxxII9rTHniUL19eSNFWeT
ySBSQu7/pRCEE/m/HcfIpPil27rTCaEMPB61wnPlrldzLu/R/KpP0MJVIsr1n/uRLuJi3OG5SEjn
NBYT8oC4UdIDPPW+oCDIVv396X+lh2WGFduUQhoXDLYvFGqyqUtwTDtAppItu6Mjs+icVSF9+oI8
IF5IOGu3jiw84n8APURdU9GB0Trs68wlyzDcl1fp03qyX2pWzp8q1DaCF6zK7/8sTpknH5Lv7NzE
4N3BYXETVeQ5B0BSilzq4DnMGa+JS+6HEvG27h+pS+7W5g288ONTegRirL3IwwLFPCHkvhEhUPIP
lxKsw2fs2nhVppuJOwziCyigRIS3sgvVz5e4dCnoVFEGYsEieuBUahaWI8tBOCijE3HqPVX66KK5
/qcjwR/S1hfdy9IQzFHdxxjqSalE3JfLFYb3DEmmQ5ezAoFvdIKSQIJRnmT3aPz/0uZ4NZ0+KpkH
Q4uL2F7a8LkH8wGjmtRkNAYL08oNtkmZDUJrz1zI94EhlmtMHxDZSAtrpdk2eopZGXG3YCnTsgVk
Oxrrn4BEHmD2DF3HRo8DS+99XZYgcpINb7UQejcb/2wgBOYExaDl8pYK7ycA1Zt33VZJKTcxCDHn
UI0N6/wCgnGFazd8LE6ygUaZ7ibUn9GGM2Jw++dDkvWRIHWspX2Dp24oDEebbssoYZC2sVC0hmKB
yf1TIfxncROcyBo8GYBaG5AENcZ7PzSzhEDC5JGt644BLGchuPVF4LnqGXqik7WmR02cSSqp5NQ4
ie5+YNnr/w91d9xt+b+xym6czASFVvFiCEn1WcwxMaJbBApZDdJhGr4126+ee4LYa0PWgwbhoLEl
2SW3Mg2j32n/c7zGgUm3djLBVSSpYDBBJD7kWYJFrkoJ1i60mo2km/DwDDzjGsP4m4Q/YY7sYRQ4
k+m0Mxnd4JYetTJpq8w6HxSihZtCCi8TbRsriI4u+a8/pYT5wfQtg+TrIoMU7EOlMUGLxw4fwXb1
RTXjsceHz13gT7YVlVQ0TbmCqPk2dExyPMaYoTRBfGnQFRESCEnchJ3bb5KaZwzCKdF/euygg1NE
G1A05fNj8+u0Xq7bGuokDBWeXHIBEPR+VkzVyD24pcp9XIvpWc60Vo4UUsKgNYyMTaAecyULE+EF
JvzCSSl4J4Se74+xOSNG8OQ7FbjoQV/+5tHp6Ryt3fOLF1hM6PgU85gZ3lYl5di2zfavcjVq/ONy
xE+RRXtMdaz/WcACbib3yZhy/ikmFTzCwvxxX1Ua3fqYPIqoRDL5x54VqHDWjgJJAyLws8j6nHKe
LF23qA5nd53ZZkeWiN7QslznndTUalen/3wN5vY2dExkAXMCiwvm/2LpioKQG9EUR2QImQEFZkZu
RxYrj3gS3undj9uTk0lf+E1DEX4CbBVytHDENp2K1935NRQCjhJRSmJrXXuEgB5m0QAlV0MKJhqb
2rJv8NuV6UGgZjtl9q2lkk6DogaRjFk7pS8r4C/dFOo+ovLvlGtg6zgYBP/3tswxgITPJlYH7Un4
cVZhCGCWonDBvyTbA4uHABoq+A/cmClsC5GqknYz0lk/lJ5sxrMdhAgHDxS5KBDbAe8JnTw0dBAo
hxs2hH7Susvhz2zgzcasXY70eB4SEphBPysrB9G3dT8YGPp8faIFsKsjrD3nXofCv51zZbyZU94m
hNyhrC9KZPXAqjXrY/9o2GJXl8q4+mJ7Xy6X4xxJd725hop1gwLFMhSMWK/JA278JZdaP0fOfFe/
yhMuaEnZ56XHrH7knYFbUZ5earDLU1g08JQWVMMeYHaD/8XKDrn4tVbdltF8bBBEclfDG7T1FLnX
nckrzFM8AyTTThf0EF9+Y+Q0UHVHbZtSFAyrzE5t0GLM34nYUMvJAjssoLyKYmdOfymwV3bsKB9k
Zxrpln8mUwQH3i8+GmoSslAQgam4OZHiH8Y2jpUEOE2bE+eXoSciXL6PYDKLoyPRqkWKgYDXmpCb
QzoKItJ9cifblAM0o/fitfeMa6RbDN/bCYn9sOBTZbVFLWnxCDWIoX+HM7oIAKCwcMsPYN5aHe+e
H6oSdbVu6z5YIZqdenBc5IxQaFW6u5gFqXLQDTcOB42MRrfhU6PBDYYIQu2ujCu/ZL5Du8RWgg3A
n8ohycIHdSlbPf3DpzP5nXPqMy10rCqnweI=
`pragma protect end_protected

