`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
o7bXVCfmobTezHsufsmCtHe70Mdnp2UYFrOanNBXg5l9oMG+MHmEdPxwIagHkpC1FekneJDtJX6D
cEVEyE8ej1IzNRd85pXVEi/P3ASGTbedhX7pDAmNQVxVbgl0MfdzCmgNl/VVp4hPLkT7AiUwuDze
pbRPPDTtAH2XTPGf6zAEkPiLnM6cjOHMFe+xp2Cdc5C/XNdVBA5/ddZTe5h9aOtNsVZnSAqwfYDN
mBJhr499HezkPW2P4vZdc8nAvTFGlx9tu0H6syIJoPQbmBWuJY+3ZITkenEMGIyGUgVAm9qCE5xd
pEWOOO99uyFr67CgqHXly1uTF5oxSGAcNAsDRw==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
tcwHFQPIwdKzYTgsk0tBkwaP5k73Euis5pt1VWlYKyGqFxKOPxFcJcYt856yNf0TQwfQvI0lWAeJ
pG24TrI1kqIUFXDt5Eu5RRp/QixwJgdxGO+MD+E4qTUnn2D/dbXhBj3VIapQ4bE+kbXUcAVpxc0B
nDOz285PZz2yooIOCnsStlD5leIIX2H+DP3zGaDJtq2ejw6MRGXu7I0/OFNkPiO2qal3nnJfXxXU
s5sffsEpn41o/lkSgFAQpI3+8h5hDHkPV9qaqGzOzoFnfYqOFMLD3hWRQC6RHZEQpptzZdjJ3/4v
WevgkyB8NnlTys+duqVJy8sHoKlhSUBP9xGhagAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
l8Z5sPyu4XvLoB1gOeEDpD40xph/bDBZ1u7S68PRUVfyL1ps+zVVVZewAJal+YZcvmGx2KwSeljY
bmKUDyZmtw==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
UyEErgJ72sK1kRSR79GI/VXYhW67eJzO1mDKyI0lO3HPsgHpAt5idxkumhezzGP1wvm6OHahOoJD
0dGSCuWGEPDtRNzS2iVqv4GivdHslRPK869r0/plijCnHAm/Z+Oa1CFhicSx39X8lOB25fWjllRY
mO3UDYULqGqV8ZIzN+WnXTNnSW3jjzsvplHw11yzh0zfTtN3R5QFg7F9xktoIqAr897hVjKkDSZo
CIktEyjxuwFVSMteM5BdXuBp3QpxlDqKWYTe1S+OT9n0Epi4Cyv9puCdT3O2XDBeOgHpkgRCgjQ2
lxQFoJ+EOuLtyiA4fgf2QqWFWQ+OtJgohM03sA==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
fJx3SMGyN+AVVV85NHzopejHi6bLTvOIK/QNe/F4mgh9xicRI+EiGNtvyceU1lZW5dj5uAUB3BLE
clSWjaVt8BeYuKB0SAIk1DV/eSjpsjaFO7UtqOxcuROWuuWfcFoxB3x/o7DMmRBKF47LdYX44W9Q
GLg/SUdTs7yhUSvCTOinOkGWxor0Y8itn7z/pLXdsAcE9S1j4nVpV4cREuUpZ6M8BjuX/szM0zEq
9SU/Pn5oVyAhTQdwgJptGvR0f/MzC4t0oiEa6d/k/k7aUI+SNwlW5SZmx5D0C4GAvMyoe0vqsOuM
6gH+gm94IhmOJJEAahiHYaLF/xYCTrJ2Tl9inA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
pzpvJnZopDOkkynJND4y5kS8rAccGvnjOx5AvKw3NxsnFblPv0N22/gmHGZKTxjqWCNWut2J/IV9
gUtIrcvsWTW7ojoHy1Btul7G3cwvhUKEw0NiodxWxi8f/oYngmpP3WxfvTnwn6QO+lP9W7Ft5Xk3
Dig78twGlbskn0/SrJo=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nujczRIP23LTK4buJGeJ+QBMj+3spdnC7DNTsGrfEEAlaYbOFXBjEBcUzbTyBwUs3Nq/ycCbMjMy
/n83yObNlQtU+m+hirGegvKpM7vfSXjEw9x7pB8/BW0Di1MhsXT+FRK0KR5Apm5q36/M8Da4953y
nzo+96C6Cx8EjQkLAlt5ABDXiTeRJi9Ji6G3R/yD0z3tgev50rKR7c/ybC/BHMTyIwRHzN2GzCNW
+Nry20wPBOlayJqFM1m7xabNeZ4jzwnaM29EzybPHIE6KlgkvwoTyGx2dXDWnofmwYZss+wxgD0X
rPUdsRl1j20MvUMahLUnUqyHHqS+n5UoWKqyDQ==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NbK014b0Ywtm90TE7zlY2Ld47TiFcuadb8W4oFnQz4dxyyLMD+gTtsq0948zX/hwn8g9IUFYLnaz
+wnacgBZo0ByMtuDEI6LLxK58Q+Vjlswz8Sixdt2eQs/psT0rYfkqlMakUR594u5Wa6233KH+tQ/
C8KUvc0aPHY2eb52qwbGADqih+6jWzN+HqTyLpkeZbLu7RD8tQlo9EeuqHn3WKiALNgL95fbaLdN
68fJgILE+b8MNSWMjfslm2crjpUnbOGsRGjXFWiCHUMQo9u4bMGHBiQsAE9kN/PCkmIIpbOblY9D
BjWkZ+sbbsZQdFMWGOXwqN8TH922wa0/yvUORw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
g3nd0CddeTP35i8EDGXRmzkh7mwslMXxYs7p82qGhMLaEspskC46/kWoX3ed3T6etvFVgssb4cYZ
9hX9Kt2U6U4UXN6ebY8zRpt/IoroQEK8gEoi8Mqor+O8V9aZfgQrXe9DHnvOMilJuiyUk3ML802+
9AactsydvXi4R+kTeng=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U3NV8rOxMfqi6oy2Ai+o790EXlbFO7YKBi2UYnmdZp1n2XfGQDjtryi893ox/TH1d8qBdofyQcSE
mAxkum+13J0DWE6K84wWe1y2Y7bjq+dXC87U2uQmjMK2IgKwSdlhcS+VCSxlykofTDTPk7k4OO5A
UiAdIpCg+cLYuLUZD47w70vqYlybgtuM74PVXGslYYjJ0Ws57cL2wskqMPf6xlIQcfOoRY1Mph0z
3e3jkiC3ki1mxCkzcu+0fmtBZQK45vThJO37jX/U/g/AUTxGRPxPPfkccxxq+/SpVI9rej0NW0SN
HabyGvt/3eEDY0E5UGRC4WMi1GJyrJHtlYCPog==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24672)
`pragma protect data_block
laCS/BCDDNSnhDK5GNheMbxU7qLVGwuc9ZDoO/w/PUZbz0IQSrZUt2pDNO/veO5NLoOu6EiZpJAX
M7l+zZx5gIct9GbeDtErluZFX2QGhln+02JF51fgtrc7qmG5o3H7bifXywUz5stxrPuWGUcVXT56
laBsTpOG9Oa3QRoiI7uTngL280aQ2N76oct0vWgpU9Z8Q61qSBKRPEOwJmmTTkJbmijSS+orbhd3
Ig5Ahec51bWPkFSuLcqjWhA28pFZVYs5CmqhUzDuoB4cCUUos8rH61uRtqsdPGvAzhqzNuvijISY
W/DKBchNnDAB4DtTdW4Un5YvNJgbduNXioGrU2aeSDBY/XQIN9iEFyCw2c4VgT3B0DIsrZMCWkMR
2LQknnG3fLYfdhicfDTiqBa7DA9ra8uxQGT7/zSSfl4n5vdMq3OApLsr9kWUNFsvGCRcH/OGbqnT
koaFwr9x2bRFfkh4ucOYz9bsEJvx6AK7LOtctAD7F7JNFrQ+tsQV733AbD3JSFFITCbo6sUen9Qa
8YOC/LdqlJRE4xYuAsrqSfDrPVpvx0j2XLr0qKwN8eO96ugcVT/WbsRTqCCnvwJrh8I8kN1DdYKR
OIjp8uXFHlfWTIg+cL7C4mD4wsfCIGum9OGW5TQ+tscRxH9TlxDO/cwoIxqyGXN3CkvhnlmGMi2u
+Z9Sl672lNMytOomj8909D2f3lNPDs5wiZBt7SBvx0i5CyuQfJeZWG2fJj68ngu3loN8ZzdhXl4p
9IVzdgdB3Gdb+HPPep24ld+UvEOaqU8hEpnzW7WnYZKN8IdH6BdV5dorqFuMG7MBGz+vsIVbS8iB
z4uu76R52ARfKsrrrRk7QPf1ytJZh3ffjF8VDGqre0HqaOgD+9OrVfbLGLzulCYWhzriLBf8oIcr
wagSK2q/HdEDo6NX/uswjWlMQeInYMOVgOjnolpJRvj9S2Ld7cJOi8Swzpsx6fQPKLLVQJ72bN+p
EpabtJ9HYF7JJKSFoUeLd7mqbuK5DPZGpadX4PpQTN1J9lCEwOCFoc0fKOh2bqnVK+AWBaO9pq4Y
r8B0+PEX9sN3pCNWegvGIe/Cgz7evE8LwHYSShcs2lh6zrgWyh5TqbPHhpLNUR54IQ+D3WhaLHwC
Hqk/IZO7D7yqKu/eIYcsBbNRUrzukhUusl8Z9cFBVk/n2R7T47wLHDhoyMJAg+H7WbN4w3DpgVgp
0nGj2hiPBMnPorkf0/XHrASC0kTewvOufjhpWUBoUwXg8Md7cZjdr+ERwjmQ/+KMkSjcjhFnHL3J
Mtxh7FIA5Q9Zc9T2fXZb6+4fgojaFF14uWOqoy20TjV45NIXY0wIkK9L1wXj3lFd/JnO1/iRfysy
NCkInBb/TR3iol+girDhogdmZKuL61x3X2JB8y/AdLoX5NafMahrPQ2X/7powoG5iSlWNKaXl35S
JGlwmLQKXFRhOTzxzmDNKUi+iS8aGRK2mrdFRWpRClCPuPYKr3YSEs42zczvt5+I541hVilPeJy5
NySA/mLqaiWJZnf1lAkGZotLRH+6Hrv0i3Wd+utZSvFa2S11mN6IJSG/k7vHgcRaZWoRGGCJ/Hvy
tzIHIOJsqPW/oqNF/zC3Jsj3WagkBXUae9N9g6Ux4X/AaHz3XgFi6Evx5Ok+RFYRQgF4Z57UyX62
G9WL128awjgDdafMIpPsrUTK1zIvSbPcLB4uLL0hPPtxoOuxLcQ27WdXjXxNDsYMAeJpe9stbQbt
pz2apJP9o5hCzzhXfQmUo0mz0tibV8ItCx3RYCU666FB6eFo/UhDgDnx8g+iScKPZlXgceydOYwH
PTIN+xkMBtCKnCMMiIpX316Awzna+ssnswZBGFUPWMmXIuBeM0vdyhxd5/RzwxvMtVmzPbivmVvS
Y5RqeyY8MbcTAYFTLCD2jujsmFL2vn0T/NQVuLxjEEW+5crm4oQ6BaOrn3bSacxvP6V4rVwd9Xrw
7b8wXpcjkWZZ5urAkFjWThUtBgDdqxSMxqCNmATPwp5XImm/gDdkJpuTP+GlenLxIIfm+zeCy+ur
5916RIDRUjjT+ZkQ0Sq+6e1XnuUv6I2wZ7+CNe2jZMyImOhPjRYfP85c41lAL2x2uNYwk3jBJME2
liScQytqkmqOIuil1Hc/WEKtHnOlWx6tilcQZPE680xp/jAmeUMVLlo7DK/ZZO8pO/dCotpFiS2C
0uG8Id7TeXrfTCkVVPwUdPQuo7WKeg4EvnMKjeHxOlYoXI1fPfioWqSjGfkIftNrVHLfzJXPBIVb
M9u6GEnEgFdcgk3vYDK+wrFFBF+RIX4+UVH7vUJ74pjko5aKdKqsfRqHn63JzP+7Oy374ll3alxc
RvwVe278uw3NcSRdeW/TnzC8XpHq7NKB5X06/Z8rvw9kLju8bizAQBxSsp7fvqDzrxKFISjEVeMj
JwD7WN3Ojd0IPuYt5YKHDArb2VwS+2J0DIFQImpSI4/kxIymj5jvSOvGNxlSi7phGmBvQz0lNKm9
l/pY6ZkKBBrwfNe2agTLCApYn8lBF7UBFw0EaQwAeted5NXNwrwwDivycc3IO+NjgTbVNcZMoMVX
dkYUMHS8NiEGU69Fwi1/C9bSHsXtc3aoZxznbX5fbxZdgpuoECfls4wjKcn8toJGvLiO2LqOgypn
0/wKNTQ77FMyduyYhNYZxn1XhleEqvwxJUqvpuBVhPFiuZr250y93QXO4JVA8Di1/R22aUfBsyr4
55n2lTrG3VnpMaizjqhxmHF7e/35q7JJFRwpc3JMoaaJY91Gz4a8nO2N1qK+J1v6FX4otnIDIKVU
iQuSaoX7loHMykc5KggXFwZHexg58JCuBJxI6Z9lH/9aVQkP53qyD14YsDWmmyO13HfxtIr6bOVR
X4LGpELTf67UVr06zEj9NeiiWyEC1aEoMJCxdGv0N3dPdoGtyrbUa2GHCNg+kHS4IB34+Kd6aq83
ECsqMpKD/ecf26oMKBU2NO1DpJ8rSQdQRqUWLAdZKdN7r8+wZ5STFnoxouiG19SdJEtnEAcXG2zu
42krHB5Iv3rt6aJovjSRMhGEWuoTJ+DOTXyXQnSy7M5zJwiNHffFy+CJ69d8bR2UhbJQZWdMLc1A
VLXgVpV4MBtCg/FAk7zILF2qZ2/6U7oPkf4Y+frrSQ+gsvR20oztPQBUzEMFQ1tE5pbPrB5kzLRn
CXHEHGW4vdOTJfOmhzlAM4R3b65AtHFGTQ4fsjKFdcUUnBU/HqdPyX1FbBIkCz1rEDdNY97cMowQ
Kzk26V4L991G58MRQzt9HbZNXpjjni+PmNA02Nyqgv72Y593TmD4nt9gOu+QVsea30fd+3qDC0Db
VALVmyhKQMvI6Xij2VNWadSikdWg25anJlwXSF21lvl0SkEYTL/xjDEvRLFTp/Qz/Y0oJz7UBYcJ
gBQYXqszqIt2VXOl6WtVdpORztfWTGa38zszy7vMxMF1lRgcc+q3FZo6M6v7DuyuaR1zNqAhjVUg
GKMN5iS6v2K+D/enQqb1zDEDM9VJu/6yt1GK/x+/gLFAMZkPGCwOtUU2Bx2ytRsnxjkOx38cLNMl
WUMmo1EnozFKeRNVv00th2rjTH0SIM8wyQ5SmImPHcNO7U8/25oUNTGxJ/z62G5Te8ae3c73KKpT
4i0DPrMKKVrDX5eNXUkoVRBgPH/fd+wy0CMnBRSaxJQE6Ragjsl8w66ZfDoX5Ej9D3X00U84g5Lo
2n+CuGGdU7szYqce+C6IsoHHa0z7KATme9Rty61h8FpIj/4z5h7P/C70Z+XVMUpYgBklXPFIG4Ni
03wYa+4xyhn22FLtmPffZcS6sXCPq8CBbqSxcpaFxLHrTHjWn/YkFR8gS29s0PMYVaGb2lmE8rJu
sIFoHdUX2mC65oP3gsoCp6P+MoDJdukKowfIOwsq8ByItkatKDdXASdwhQylAYbRWb7j1LzwQ6qU
rDZMIZYTz8+4kw6AfKP0saQStaA6qek/bZ1wJXnH8orlqS4Bnh5KT+hKl3O2E1MQm3/dl40+QeOO
tghS/Y7oDAoQ773O/+jjLfdynbYSE/AfjlK6NZSSvJHnGf0fVc3GnZX3eCcgwAFy7kbCexwrcVc0
zqMKtvej3Le7um0rrqtT7k9cH42dIp9D+R3C+cZx3IMPKbqFc4KCHPxzsU53esk7poZOXkRGrAtn
cs39cfji6rnnvttRGqHIuVPdNdwz0B1DNnjgw3Ezn/PzUUewHwWiKvzhHFsyGURQ6oWMXLKPXNIT
6OMaq3ocUn1urpGUhg37xjR0nKCZbDw3J5NrMfyEFQXOUzAKdO3KEcKYpOHJTvcovS3xmHnQ5BIO
awEfU3nYA1n5mmcRC9iXB2Afs2J69+O4wvstcPRvYg57g9LEi/FCds7oEHI4k9xW9feL+sgNChtq
LwwPiku+e/PDvygWDyRbKo0ZyWUV42E8bvD7Usio/dFDnpqkLWSb/S8F1idxLv3nz2ZZO6dO6hah
xX8Vi3aPVqwWmxl+/RSpeOTkEwWaKK2ybXYDAcJXtWQqOa5TdEc1aWW9Ka5IaLvprEzb+0O3J8ie
sjXcfdcv8Ac5Y6z1myzeSgsomzqztfnp7BQq0VExdUgDq5Pu9Ut4z1HNPz+z66oKcuowYhAVD8uv
4ZBBczgvoVR6X6cHbkBXZ42fd75u631VfwgHAhEUqW5ukiPyNVZfQj2aGMWdPCQxGRLTUgQeBAxb
ZbrgU6Uv8fxyR2HmPQ9f5Fnd1Lh3YohgEZvSCCyS/vlCxrWUcMeoT6WlCWOQktP1u5bWyRyHB/Hn
huee6rzqmMc7iHapqgWmwRLWgctOKOziVqr9P5T8O4LcxM9kR4dLgcxGuAnI0AlT2HDJejDm99W0
Kl926Z1JtVuDQC3+GITFmTnQinwHgFEEFfv9Edq7jYuvbc/jN4aaKQShirBn0Mz1YYQfluJhb3Bo
kapOT6P02u2vV5uCe+Ak6sZymGC98NqxOK07e6evt/ft5LXlLy5ATsUil4g7FSt1amgnoJK25dLo
5KDhk4g47T9JeqNkJld0AeXgBR4CRfZyjd+VqwycdcMZp1F87d7xAD9EkRJ7HlQaB83iZTwRLnet
3Fvpew+4inb3GYPCbaBJrAD79QRtlattw5ndrrOcyKZbCx39RJUg5qqqnsfeZkJtj9lQzRVOOu9S
OmJpvVfrKqwVcPkdmvKWFIxvdyr2qe7fnbkt0ILcbLhrBlgbi9AH4n49ATZwJzC8PHZX4PwNxMQz
SjmsbKySr2GP7bBiSFnHri2WAWcD04EPcy5xemfZUtCLGdfziI+JbCEA2MK5teHnWH+4PTa8/8sy
3LxX+h6gYsddbgTU5lq3gjXebaMUPyE3V2I2EyFmkeWNM51KT0K4AzZWqu/ZscQXEPCB1ZOtHuqg
AqweqmyTEGoTBWhn8Fh1RaS+0iDntzbVoSI790aBEKim3JFrLiBN7XHJaAMlvGJCfa91HkLpHRXx
u1mG6UXtAki317nzMFMqSg9vY0vbIk/7fn8yczCLknQ385eFNvzi9VdgiRQN84V7IfMc1b+t0C20
EoUJtv7M8ZmkmfzENl9ZSVzsbIgtl51C+K+WD4MbHOhAiFSyeKqQO0nfbz3KE2BA4g9YwqM5bmq9
SziP2vhldkOKXXg3u8wmvev6lzrAvJE85uitPPFPIuzna4jc2q0PAQCB4kZjkq0cU4Pr2y4iWyIL
m+FpsOfK4LFUd9GYrnqdG+ATdbKzOTKlHFe54wbSAvk03wkOpGBRk3AzUESL+2CWggQgIb8w/WGV
oQm8Nf58EaKQW6JlGWR8bo4rEoDJlEN/m/Z7alDcQ6Ul1cMspK3uKSXHulS/So55EUVPQILLimHy
jvyzue4AI84yf9B0BO32iEB5g0ZZbAc0asMFAWTo8ah5ddSxBQenfuGEr70zAdv4rsmYYEwmLSfs
24OU5drxiIA7xnIR8e0DV3kx1rSPnJkQ43Rb1LMEqoUDoY5i3/LSghuxfUgBHvhIXWPGIjc7u9LW
1tP0Tc8Qq2UDQ//1/Y/6pYMFSJpJs8nIA8aS5I/mxXgr4sPV+Ro37bdOHvnzdrD+4X1xoqa+nkR8
SIp+2oV5j9iwzAJCs8jS5j7xvnJhmj+DD8CihqJyXsS0L8OIyj38iKY9exgeaABi3ffpyXYohVCD
FJ3XwraeTlbPasd2T/bntLkKyYutk7/tHGJDdUU4CObFXfKArigfbl7dAhikRxTm8XwpyHZqh0or
yJgL4AkHqUziOmb49XcvXf2cUYb8HQUqEh2d2XyDpb3ZHuMP/1c0adSVtfaVgRlPSHJuxSoMVe3q
DKA6scQUDwEG8oavEqzUu8Ijkl9ZK6Bq2JeHI2E7haPuBI0LiQd1l8O1VVXgyspeDt3Y16CAfI8g
MzpiAZXmZVQE2NK2pt0Hffm/AAlhBDtKtCedlhWtm04bcN2oozphxxGSJ66AcQha9q8nSJ2SC/ut
Ex9PmloBPzzB8Bk6NjY2EPRf6iEXWcUwCStzaLnAImQBNndO9TsqAXtqozSeU2TUCcafue62Gtmk
cV6zFXD2IGREkg/BGFwL5WK9VI/8GlVxjBdauNaefUfFLR2WXOHYj1jBLz21LPclGzchoLIdt0i8
3bJjoARbjThO6DUB7lLDNExj/iiUz6F8H3Gud9Lisk0WZdJifbEm3yJ4GocbQRgu1hOhnfWAxylH
MwqPdWXyjd80bnTAx4AWboA7FzEPtNj907zc0cSroebRYU0nUTMH8WUQfYmBqPTSHnf27yHlgyL6
6VEyrsmiNQGu6tJTdemZmQWdt4DvCPcjWC0q91X//Zapwypb2LOK2OYnZqtKELqgyJMSkv5zwwCG
zNCmetMHIVIVeUGuziblGnmGPT2omwsFQzB0iVSD+RNWRU3tXmIv7b2EMA8ta7e0VEIq5qJ1fcmJ
Lbsi9RjdnoY13y2K7Z9GhD5DpMuTk+wg/B/4ZDALBAC9+xMO5obf741P/IXJ5g7RowK4DxIQQeBm
+oHUblKWKkky7izVY4F7LXMfLTOlX8zj/5ndD5wYviCUZ2+hKtcsWzBUQjR4FMIfMc7DavES6QQr
S6Nw9rD6hvPTfDQwzr22BuU7/az+Wgn89xe+i0RAm5Cp+WiyhXMbL5h4w+2Ex502MAVVF/Eiv7HZ
nUjXoEQCLL0C5xwr8HlWCTzhHbRAt+eKt47zSJP7P870v5Sd7Cdj3Ykr5limM9w2+qq8Tsu4NH6b
85oEODQ3XJgAf8mrXurcXG2ge1QEFgciZ4dMPF1EC4d9c+YB4qY0f+F7I6qOseTCI5gHLdZRCTVm
xC9oStD0iruvB9e2+0LL+VxRam03TNfjbZCvatJmz8hGUjKQanuQoaxC4xTjnaUbx4dVWnu2pKOu
lZ/Ai0SZgTUqdOhcv9H8wLqdLawwA6c9N+t+GEti5vl4wjzUAAFhdwLuwL4DA4Hau4RLGKQEHUsB
U5+1628G4DxkKzuBbynpTcf/76V5RQaOZLQUIkJ1vBfeHMIZabP6OyQ++FzyZMGu7zEjyEe1dvPv
9KgZfQCtUZN6yJFYa9a6Sj1CNjtp96FJjdSyB75dM1QUa9LFv1L8h6UqufjuNKKaNoyRftmDl6hg
V3h8x6nuW7AdRZvMkwcex1GxmW74q2auqbFyVI0MAKBujxGBANveQhur+xz8BkVkiCrx5TFgpq8F
+TwsfOaURwi9DAypyKz9JKNauOtCYEiVZ+9LfhVRDiCGkqwrpe6vTzDrbxQzclT7Li5CEVjqlU5D
X7I+Yllc/BQGJpYuwlJTajifG+vjqkgf5uhS3LL48sIKxFvZ3Xhhju84KWxYrkMYrIL4K9Aoguhz
Q8pJo4JsXiQgw4LLIejyph8byK+2KLC/tCs/P3EJf0wCPiQj1k3KLXqI1Dp+sop01pLgGGqBzCsb
QUigN/nNXVYSPw9dCwmeaqFbLRVLt243pVrG/6ixw4KaSUPbSDkqyY+fuLDyGzGxiq3Cp9CWCJ6R
GbNpPM+MvyKKuPlTeHXSAvh3h/mNDca4OK+AxTBSTJUr6up67JKZayNi8X+Fdxt9bhmZEBXlpCqi
SeWNiZ9HBsHEqXOTfjiK+BGR3oEdRjAfBWLiDQ1qebXOiS6JZtmWjow0thR7W7YJ0hcvBa7WOtpl
TkNT3DaBd5z0IdrOw5fTs9HzI3fE5TUY1zWJ4XOTO+WkHSnNpHAsObkmCVxfbgys8UJQ2O7UVIGl
SUs4TMh+EEXo6yXxNBwVbf2QjKJryOjrG+P8s8TanHWfXWQvGe5JbI6E8yWWGlu06a0BAw2OYZY1
zxZbS8+esN3N+gL+6PGycXXPYTXnu+23DC5mop07M6FuRST1YpIybJHppbfwPVp48ND2Wo4M8HDg
87jRQcI/ttzV99g4SJsP84wP6lCWmEmIpk82gXxuoNgBvnw3gCyJVt1tD0i+15kjCriF84e7MVIO
/kkX1pgfou0ClYjtu4SQs5NinZ+lYuTNBnIUZUGHe45DamsiIwJNDDl4pcyoV8Ymvg3SCYvN9ZVb
Af4Y7CdDoOz9QWHSDDXUuJlqoeC6ZlWphY4ik+A4/VzIVXrKzjgxUWmy5qcOp9mZXD4FeBUSaR/y
8+WRTrOqElHSDLLf/6l0scdZdc0lRTdgnYdM9YSngEhFKI3U24MVIA8NvUCJtxrGNIRZcCe1xqj8
JCbbVGZSv0smzbqdOw9H2o4DGHR0WFUD0IUcvDEqEVjEZkQ2nqCq37G3MRJ0UxJ2EbUiwTQTxYNu
I+DhHA/86dUrJvu3sF+UqUS1tqQNfvEguS2LC0L5TZSkmY8jgG0FYnpJxj4E+dv6xXwmJgb42pyj
JHVavYJjOulUJzs8P2b0pYo2Ah0kKAjL2pYFUKutp3Ma7TgT6vpX1z0LR2Kw8WmgHZa7bj/Pring
0WfQz5XwMnQqALsThft6Si1PCMYTENm/lB3pgZmGmiYPQxQkk7L9wHJCnz+x/ClyrQsi/cEtu1AA
ZMMsq+wPZSPOwAvRFRIAzO6M0YdMYtMCk2R+9svaFgX1YVoOHiIGykqd5odjsUwA23B9ClFJGSYb
V/neRWWOghLegQS/XJKqXOFee2cNf0sS8q+/2Zxfyk5EPEyddB1aFBWHDTa9JBjtiFSUi7OFrtYv
RDG97Fn27d1DCrS34DbfWJP3U3pQV4bKLHDBd0/J2cmevJpQVcKVIwrfdthAWnLOg+EFafPwWkaW
91iXKyfLZBCg/VmJeaedfHAHEOxqgGJ1Xte9cvhyRtOYFNB8cldPwGVGJ++B40MptBcwXtFbRXgj
sfahDYONwDdfawl/bdFPfVMX861FXSdBj7HPp+8eYdvsZAPcGNAVAOG/gYzhPdOc9DnlFxZjenF4
GkaRx97cZvr/ySRB86qT2sKado1JdToAQuYUgNP6sK6ALgWt7fr3FVBufh2oDedht7Ui6fEfx8nJ
3pOStlhO1HGCUIgdSkUG+kpaQg1p97ht98HpfI8n16N+t8jClmGqki4cUO6OIIBzZCwPrPtbnjOj
xVgDD6chn+/Hhcvpe2ewVospASKmc7YQAZ2WdelWL326jIVtNgOyac156IF+Ao9Vu5ArqY972+As
djLKfoOMpN5FZhMny/Ks2LSwuW7jBa2sYses6PrIKsvUa+H3fiWaNQ+Bz9VDn6bNTnf34AQpHLZ/
H1iG/bXMS1yNzOA+n24kjDdPXGfalECpylLGSnhM62iiF73KSFJH9ZMvJ+SSt9m6AICsOvERR5x4
Fb8+MepOgSWcaY20NwsSmhCuAK3hh7zvqkRpONRlTtHl8+h9vwrKmkmKSxuA19BsEVcFZwE+Heww
ZoBYvZlTEvDnvW5F9EQKYmvcJXD3lheTBXpaYTSDyy/gVGj7eTfXQHPGKstf/LsyUkNhYnHrFFnd
oIRbsNoQ/gBi8SbjcToCEsW8aI+HA8XOWD7cH8eiPYMC+P87X82kXYmyMnPhHUq+UNy0BIk7smH/
7OFgSj+TdlapmFVusLkKhKrLYwwL2B7fa/DfoFjpL0Bo7WGmUMETGrYCj8Qn5pYq1hadgeYn15Vf
406hwd6GVkLSqy9t4CBoQ61kUO2Ya8XhdEuoMg8soOdY7gNlxuyPR7sI4trvAY95CL/J2KUMWj4W
kCbjbErHB15DQzhGNxkHSWxnmHtq67mZlVqWtzdEY0IuJkw/84+IcHIt06pmf/CX16WanxRfj3KU
TFQRPrTTt6gTfs0lJNME9At4qjQVhUSzVcP96wTW7lQCsJKoWR0kbQGbPnIIkBHxmhrZwXU+/YJi
rrplys9eJAU9ygjSbVpN10djwPKl660GKkxWewN52VpefY/xlXGKj3jOrmNlCMJEHOin6fUTocAk
AvKWEv+Yvdej9fkf7f5gO8f9b2xmzvNkJgwzLG613WSwdJGGW0TWLxLo33+UWfpmeu1p08tzboZq
9M+UQSavUzCCccgY6FYzJuhOTntrHoOtfziTC7mJMNiv0u9iJ1ixzdUwB+ZaGF91x8q208IJbYun
/mo5DYs/Js1v87lziLbJNEkilEZyl1fvs958ewm5ZeRvQCQlpCl3NyLDVY3UQklm1xhJJvwEP0Cf
HQo17OeFOCzEH1KzXa/aAqw03msKF3N47mX0RCX6R1IMdNPEwf3IhTcs9Y/Ens5VyVlhY4eyJvA+
IlDjNGbqiUvle7/yNruRdw0vzOcnA2ErQ447/g9J+O7Ckt8BxstlvvdWgB1UdPqHgwGHu6owjfW2
4+A+CE5gVWKmie3pwbMihb5bE2Koivb7HRgQhNkvMtUf3rOuW71gEyKr3cRy3OJ56Dwk2YGte6co
svcJJpCaV+S2N+LV8/ibuPZTyNcQkmmC6ZwI09yGcvqoEgZrpACqW1akZQ5Hqf9P3u4v52POA8IW
DuOmKnGuVFWwBnkCRwKIYNwCZCvg9yAz7P0q3++RpbLrxhYt3Jdwcx992mx6KW7hp4ZV1Nes4vga
XmhwNWcqXna7wYs0EqidOeR5vcHE+dfL4HiGI7cenwPHVSMOEyGTR8HRK/UoaHE/vIGOwUqH11di
YWHS/OuD8tQx5bEBaJfs0Cj6BlHWDbNNt5SC0at2mVfMRHLWB2no2zr0IQKZ9p3jHT6tEroOVsaz
J7e6u9ht6fpIKS/d0whPahSy5OiCFHvPV3TNF/EnFYk02bm24Jl1ofc6FPnnKHdMx4TAGM5dSTTB
A9lM3Sb6PQTh9++h32ndYX9WZE/9L1YFXvZFFYYuMx2hZzp37wBuADFpJZVwUczKF8UfePJs2w7F
w0Q2njBWQue0IJU8K5rNxwMfxsFtR0Qz9cKg3Qa7EPr7cYuX3qDgmaWPZQJMDu1DDE9ULvcQfuBV
+W9voN42Vm7SH3viBeAY9Wb0wni+SUpV7zi4jMstRrTd5CpqPS+11POWxGrUYKmC9Z8b1YDw+wbA
FKSCZc7Z6TgdO+FHsl18zwZKq8EClqZjZbAjDkWHd/AjyfvzJsyt5WY95Nt2oXdxfG3MwUgjnjNB
UroSg6Lk001PW+lhOxWwpd5QgdniD9H8EpmRljEKUPrvOLnpErd0xv9ShDXwIB7N6UerPr3GNiYG
oiNvBrojvvkR8zysKTkOsARfrldq2Nym0zr7e099CloA2s+4f6wOb0OIqqN/0bnbEASs9qe/PE6y
SJF1DoE9SAm1KqGCkSlip6jHjiAeOqpkdJa7NJj6YUoxL3R+iJ0mG1BrVH6SXFvG+T8k0wd5lkKF
h1OXf9yL4LjmbFcUrtlI1GTM3pWZztxNy8+9sAarM3bvAp7pSFlxHgwM9lIQSDrbATZTwu/gYa3D
m6XJVUS0mzZ8Lgrhn35trkLXZ/8Gig2ZKJIrlT/uJWPjK9L1BGyFhXIFL+Q4/S9l3HK1Gu2Jb3JH
K0u1FYEkgziQ5jaMqgCvPGFZy49cBj20zkRU12Moa5NQt5licF9ToLGJj3Ah7bNAR5RW5tMNM4Ug
FZmoPPsYzesfYjkBvITGqARHoCvFK2wtZNMeTRHMHq3J898qDIw39TjEDqGMPdfx1vfn/uHR6Gde
nfe8ljwo94oa0J8uMWdvDUEo43l2YbxWiMBdVY7xhWohMELF4C9e1x3dmXKUFBvkTlfRQTUEW6QM
KEbgr73ZZNEfT+oa7iKg3/TjqYqHVscSWyZ7pPk33VkaNgzvOP+sfN7U/XT6e+f9vZ83IVlHezko
ZY0rCi5H3e23qN8DfBCmWvZzxL0fu9wA6G6pVp1jnc+JA7STNHXyPan2UTzNy+x0DDINqVqZGc1R
AgFVzdto3TqdLlv+Un6QdHUheDfoFpqh7o4giHLQ8w9XjPXkMNYLj5OONm8fK7ETMbyFKGo/ipPN
CGtLWrADcxd5MAtO45rDIB8tDZPmoNfhzoRejB1tnUjm/4UUPD1HgXeceAYwERhiune2SBFv3/OD
4v1MDNpHBOVzDCVKE0wlNX+zqXmwWJBb+FZxzWHn7D+IJgiqENXhddjSpAgveWidoMECOoGbAexo
vaBqln+xaKPrUS9OezaAzN+DQzNnEGdRhGPnQ+98e6g3NDYCYaxKstzAwckNJ0Co8NKPZqIjRNoU
h5XucSKpBe3ncqZC9uidC/N0OfVx0HWarFhY/4F1WAmdPoYbevHEVciFet0HJZb/i9KhtLXXXJcB
oK0wLpfjZygZgeNuneQKCbwNtLGg5cX7rYAzYn4xfKPbNe/fJq1UKCoeSxLel3GddVxjy/yxjhaQ
14OvPZdZhmWZy1Q4EgTz3gvBHbHbo9knSKdzilKsyp7AJAMasvpFOKk+68tt49ic46QxN/h31Oqf
diqX6ESGifRbondhhR9QYXHOGXggyWzw5s68oXeACEJV0KsgkRAzeuoSjHXb02sEptCTjDMBfTmO
eFnkuw0/B8uhwb4x2nWz4mBmKfIASYLMGQDh0d06zKsEk5nVbFirmH4J0wU1zo0PD1TRwSDNDK4h
LdHK/NwP+qBuhuFTYcWBWCIvgVkYOCmwnuqIkLuKgvvFSLVE6rOWKGmbCroh6ljKWnxkgeaFIB5Z
4SSPU1doO1eFwI2o8qag2HDsJOaB512eRuGBgMN4GXlgrevyD4rK6fi26xaQvAasn7a4nkvv7rdp
N68Q7zQwHaSjLrVJ5C+wisfmxLp3fztSphDez9sIwaBVizfoRufL+pI7ekO/8xckVtjlJbsrQVM+
IoQrGw2c1ToSCzxu5Rp2tf4fI4Q6zifS96ifmhEj3mZCD9f9zLNz/FMFZVWgJnMvwmc+vtqQBjTh
85NferdZ264LkNtx+Fz2pSZ+/OwmTqsZupB6clF5h9IgRj9/+0AqwMC9oRqsq+BG+5/f6bcDMxZ6
0agGcd0fnnUOz4sHzPY7opieJ0qTF0JN4EF0S5rR6mDC6v4ZaVmSDCawEqVME8c03S/Fnc+1VPj/
4fUKSiY5Pi+cG4JZPFS05TZzWycxysX6G2rDvATuVnljQggNFvS1GXesUc3Sh9baSl2ID7ONRuYz
Oojc2KsBg+oWeyJbOt0BW21VyTuzrwWngl4MWi1lJtd+g9drEKRKEGoF0PF0/ZMfkSr4ausdVLvo
DL5UAEmR8GjwwYZ+2udeziySCHdqzHWGiraIIzGkq9r85w/P7bFYT3BRiVVVq7YWtl9vuz3EscAN
bXorGNFiT6IAlO04NrWVYV9EE0v7/FFywePhXwbWXIf0F8HOyjCGCr/jG4Nb+Qwca0Ndd6IV4cu5
3X6n82j1zDDAs49O0NujYnKvn5qn827ypHWo765ZAS432D1rDzD/jsP6kODpQnNpt4E2ND+s7GJU
0rcLi63khSdOhpBoDNJltU+C2tVE/27chNivcgGL+XXEB42zLX1PhvZOG1X9R7t7/QmDLuKn8/FY
+6pnfYbo/+xh0Xt1lji3o1QcutIKJsEg6DLUdPEUXDXzA4T+ZAHfrm59Tyu4UM05uZ0DW0EeaV8E
Y0QzwMXNqIM8YNntDLLjgxwwhQi232U3fwskCJs9uJpNBk37YF4aRxNqnOd3mEMnkNRObT235YSx
R/BQcex16WjEPBf5639lJ92l+iBn/Ea/26YuzNvijfA1BzW+1PqDOOF7YkQm4U6Qw7psgNmYCuhr
m/Z5sIuXgJaSxdDvMBecfYU4Hjr6kt9Yy2AaCg3nle1RNxZu/3Y0OfIvkKKYga7WNZMDGhbG0iAO
xfNV5WU+zqN+TrKESGBR31kL9Qfx8hscZGRN4AbF8d0+ozupwF+3bwZFc6Dr0WWkyLyK2jkYlPQE
0NgP0nTfa7hCcm4eneU3duUlD7he3E8o4xs5po5DptNEOXThzz7kcEYCxHvU73NS+NVXV/5RHUxm
vFwdUd9lrB1w//I8GFD2i+yE4/2Dz/7BntD6pcRMwBsvwfZOHJKBdbpOpE9HfQMePKUqdja/GDCy
r9m0UOkYO9YwL/lGbdCPzplBuQEZQ9Q5k81Q3YQe5B1KA5vgQlWB8fKxSASocihTafOcs3kXo/hU
2zCjVgD4JTSa+PEK7nlBrmn8DBUdPsCa0gVWl2bPgG/ysYOZczS59499yTS4lU/Tdp6KydyGL2h4
+VrVCKIOqpBQRs119CBtTz30Z5mGkNfHNhGlRN3u4t6Yv4AJV/udmG0lq/obpTH8qEFX11qbD4Kq
tQkyokOWg+EdrXC+seVR05TSk5wLc9jbUpvs0cMJZBRTWVGkVIgHB9SI6HeHt3hgEXCkzwPigp60
S0UjaeNoXxMPQgerna4W+L2E8Ef8EpnooWJA0KOjgBxBTlrI7VxLjp8gHBXyvnPr9BKw4OoNp1yC
Nwmh6WSeAYpuhCFlQ2Qh+WkOhSdKsL88SpTSrcjTzpQo4u6hE/5yRpsE9InmkXSBM2iu6dzOn7eu
Ot9N8Pitn9UyXn98DbxcikIvxzMgSf2RMda/hj9NhJocGF0bT5yw9U5zbyuFmS+CgXRuY8kKMQFZ
1/Nm/w0QfdgMoJkJYz/41mmHxdua5pPdkQxlXCvKRSM80e2twOTSoCaShy/XZBqvO62mYL/Hq1Kc
xfhGuUt9R9JadWqcf5gTdcgpcH51+6wS1ppbloj1ZL84/+XG+Ns6KeRQwneFLZldUCq7f+sy48AA
Wq0BSSn0ePcJuGLO1FxJHRdqZSsB79RUNkgai5TfaE+ItLLplc3DXgF5X8cTsKP1cGlE8Ii3h2Wk
2azzi+gcKvjnpVWa3S8n0xaUuzKLIP4glEUDBWdGLk2z6s24cm1e3Fnq+aNUw6xD+MrxOAiTdw/m
TVpUDTfEjvoMTH4xX1qr9PHYyWOB1Mv7bij5EsLJKHJrzI4i7RINnepZ2lgFfuxkz1gF8lQtHp8J
s7uISygd2CBXkhIlrB1nKfZ5lJCv5xCoAUQhYRoXLRt8bz5SwV7QOOznq6nhE0GkBqXMwUUP8i3I
Kujtns9JwaMMZvn9GJVacZBKg5mxsahNs0Lhkbtoc0n0NVqh4Ic1py+p5cIacYw5P0Mt6yTe10Cl
rNB6BWMUsFM+jjPdYwjZNJ06XISFIVa0utvdC3SfLQhr+iw9u+TIuyIAcLzUX9FXFhdlVJP++T23
zxiSNzau3UrwjqPUiSg+BZx0XmBGw94jFBh+MGAap4tSo1DY37IltWjeXsjRd9F1l/s6K2HQV4Zi
ogPYRLVyhR9G35/Sxlq/oc3IOijRNpWXCMMnHtlmPLNLfJqDxT+OjNSFOECZDQz1SFJeCKcyG+v0
wqONRZVMkKOy1ocJZlvBCDXmkYJgOGKNiO3d3kgCkBFT4fGIm28Zbm13i/3hTd+YmEbBERFbZ/Y9
T5HjynTrdBURisfIyD5Oq8chZ4sguZO1dyLuCLvp5LEcxvc9HtcMUsZlZPVD8mWOwclwmwGR2YwW
QDAq0VB+etJDr7TRktwzhRv79B6ybe+bSL6xZXV53NuUS7kKJSPfIC0AP53SyqVXpo4JSRj+pTNx
UPtG89c+kNuMWqknpv9kbnxMQ5puQdwDByh0/ZWANccFaGwrgWqXTrzmIPH5LPNvxAY/AmvlxdkQ
yeRjubmhmbRczQ+MHwAh+q8E35c+O2PONCw17hd87b3wdkqRMTzUnkn5hGoXvxQjvxx7TccdzRdV
zx+dRfxeI0KTsG9JpQa2wBfl7oyATfWoQmnx1KXM6MJrImwt8u0LW40gPjhgJT9VMS4eXODjxhN8
3ByAL+tHJXxqgLrNx9QIxzrdb9r9suETKSGq91FfwRlM8q9XBSRFShKUhHGJGOXcWrKkaTdwAosE
vNLcdDanDY/U3rYbpqOA/n5rcRZAmcM9lnXphUxD8RIcvIaIvY5B7uhWaX2R3Na/J0IzVodgL8f3
UzVxwQ+ebEYDD/yKLQSSIV/eYagwM5zGUx3jGweRScTrRWTdEbYM7/V1DtQnnLInSlZ3U7nlITLP
N/PgeApJ1GIqjbWOjM0a4l7NapM7UTmvLiYcHhaeKzEx8vhd5Wb+U9PpUNrA+WQ/GeYxCgONZZt8
w1ca78iK5GSLgV/F+S3Tu/ib+wlPdcatNGpbeDV9WEBRuH7r7dEmaBeFdkMFpvohZ8J5WIg5E1su
4vdm2u9+vGcbMtgetZgnzDuCJpWy5U1VhzrGja3aoJiltN2U2JFSvqHptqaVkWKM2q6vy7NErJOc
4+VVNlGe1xE9VC8jBGKxYLgkzE9r15lJb2bqE7aU9vod3+P/egfp2YiXGZ2wt9yMdI/Aw6Wyuvwh
kfJxp0owGPsNhV3mMX69ze9yzWli40zDAU0fS0LD2I0UJxYduHnwBOug7mNhYjV9oRDE52qICt4N
1DNTjYl5YabgQHhX+kqz9M1plip6FebGNe3e5Q1ZrjEiRAwKuI31kweFCuoP/oSTj5RpxR28gHSd
uCnEvnstXc3NmhYVGhCJCfK18zspvzhQxFfAS/NaR2xTQMuW5nkDet6kQodUODZoJ9uJKMzJMo5M
lh0V3k4Z83sm19c4RoOS0zFIF/UxeXVhgPhhw1xF7ZRNeZtGSE588MPMQx/e0QocWHw+9mICkXjr
pSRErm4DnmN82ssp+8+v2LdxWb7OL8xiJXQvmepdiXb7CSOmfVHc8elwn4aegVd/Dv3R+XIW+SPW
6LmASqIJ9l+JFHQdc0jr2FmnJFvGFNewERFeqoUx9NvAG0Nl8kkgl18tJcxXZp7L37DZKAJBW4dM
PfiHlgi1KyLjKwHmw2AMFwaL22ruE9igia+R1j4X5i1dtn9dH4GCU56UgUfJxd8HBj26aswzvdQV
xnxZ3+D5QXKB7ibPPhQNX2Wq32d1aT7AxjsRgXPx+XUrF9VJvzhiFy4QmagZPcr6lLfZcqaheOzq
h56VKpC+iLYRmbcaYpxweGmMEP6XdD9j/1QUEJmzB/zw94xOMXMu8q88ISPnaQosTe/98y2Ti4Xa
5jH0DAvo/pcyLjxHtegbLC8Z7fJeepDI4VkA6GHFPHeXaRkPfqtIPobAwWE93rnj2JBZcJ+74w6m
s+6jO0WaZPsCJaZYDugJBfsZPV4NjjIxf0vwSpGKOFfumYuPZ1w6mUyG6/XstOPGw3r2xlVG5ifd
BOjs0j6gzwdQQpS/hIzE0KCidsMSMcC84elPBJvgQku76JxNADmtSSvi8+EtIHUag5+De5z37bjZ
GGa/RiOf2/NgMUOJg0R6AsHbXwG/DppXZkWdO1quqYQCT/7yz1xGw4ENVnLdtNFxYhNeTRIQWBGp
KUqagqA3ziBerLJuPsYxB2C6kUQGVOoP6+Or/NQp94tbORLzJd7cpRh0yQSCNMkXJiWFZ/XdtrAj
YFfRKb9obRKy8TWr5Yjebu+Hd+GX3zNLbMCd7JWfoe0sflItHwQGYWN/D60NOtQi+Qfo06pvlhoA
nvXbFLxoQgF4dYN18E2ktRX32lwdxhRuOc1IP84rdFyHhCyMHuYnNs/YsrB0UGUFvzMT0X/bbRUu
S+6ESq0NavGhBITBbyhAI2I38xN+LRCyBHMjNsLBfWZWZ8FMTuQF8dp8q5/oMHvCX5qU8yQswtQd
Og0TWeqN0viEd20xYEs2PbSudedfSYnTpmsVhcz/dL+SzPeAyqPVNjrCxrYpsCPQIJtWNA1OzWjn
i+owkDUy1FHbDDG+jI/54oQ6SitxL5JIbJ9emNnokK+hjqezl5B9wDD7PulzWM/xbM7sdPTsor7q
YsbWJLhKbil45FHJaLtCPajd6UfySBDpNaTANZ81Xh+udhdz7czSCG0a1D/I3vx+oPxQrhRGIs/c
jlR8/IIlGBaRlKMbNx9VUvEee1F7NE2/uDPMEq0pJevfbK071ollNAja8ZkNI7Rriw+ofCyI6wVk
ByBMPVGTiM6XIjJzCfa9yyolxAgURYAHKof+WYsxH+c+tOl1OVMfUCXk2OyVFbPC3b0fozWxzMKt
jmh6GPrSY8In6vpVELCM/FQyq/oyVQM098CSif4QfBdUVfUDPFLWUcm/mazjOOV1fG48mexntKoj
v6o39EoAJ+3OpERWXY1RiGuKDQtvGDfqxj4o4bgnlJIPLTOOvvWHm6vQySqLmjsEvz+fat2yDh7r
T7tTzCxeQ6Ktf8/HYe9ykLKiZJ+6KvGvTvsV9qtl6Wd7vXUQ/AzoClt6P1GdSPpRGJ4Re6o4o2PT
2VTk9S2+405HeXnec+hWus3a51dMDJkRRYpR3iX9DTYercC+YacIvquSWSSTpUiqPWk1lgDnUkoM
l41oDA6SRDyWooMEhKrOm7BDcm0Oie28lhk7bJ0Ug1SfA51tZQkkC18p/X0BanGE3qjRTnbAkNfE
Cm+Zbka0bdmUeWiy3hiCr6ct5N8YT5RGQCs0o0PxGYYiUwaQaBokGkPtnoNfgwl0wAmvN50Kuryu
kxqIofOHaGDGcOFXhR661DyH3/dcaaMKBdupTJja02VR+LdL/d5K9P58RiUXPxQcXRJISM8pL56o
8k4kOOMVO3kEXrRDaDbY/8aqQObqEo+WtdQJwNplZqHYNjgj6KKSnihaYxWclHDTfC8eJwxP1eQ2
vwtY8IbGgGfPsNfx2a/r/cyVvMj0KClf25W1vhEwXMOYaGApXi8MLTj+RVWYDK9EBpeRdiiyBWKk
v3Ip44KqnDTnBMd3PyYaQi9F5aQC5eoVx2a0Tooc1sGVksnGH+/h7x81db/pZnSELgTuJ7EMJQMh
Nhd531pa3juk+/16BtAsvGIS6S7qYX82JMCvUMRyrsjfXjGdYp9oB2EC5wHsSeX/i9sNoPAt2Yiu
GIWdZEZQc6/GadyV5uHr5Alw0RWVTBCQCpOpetbJjNiD0qvtNjV51WUOJIMj+q5tiJAI0xJMg9pG
0QF6XjXMUuGMgc/yjAzVFFrDweiTn0E8YsjsDYrkvYaejeOxBnx01iPGM3wp973gaUmU/6nhEiC4
Tu+VfjxKBbCckcXX7vTEq/Ti4Ku3RIOrOs+pn3nEbvvSliiTADd3f8E49YiMsCaJw0gCtL6NqfyJ
5Z/bd9W8dQbyqJr1WzMRHoU7qMvoJTuwvXKa8xJKwMlZXEtmtFdDI8hVDpcVR/fnJEKBe/0gEEe/
r3Q7evNCT5bJK1R3jBokVWOdf23bG+x7ZamsrSxzvm6F7apsCbkTEkl+f1BY9Z0o3KVgi3Z4Z4k0
u7l5JwrPoKI0B3Zyao2XjlH/Gyys1eYAigo2+3EL0XRNZ/lJzCJAxlGCEx1Z8+WpoRKra/FzT6+U
/gQpmV1UQgwouu88S/dE/gbjzKsq54lsGWRVfCVC+j/xE09M4RD4AhJye3Z2blYLjN3cG3FGqyg3
lvEuAkl99ro6s2qm/+v/hYVTBr/ZkmSznUBx5QJ10BfmiIgYv8QKXcO42kgcPXgrbH+hS/9CrC1z
UZi9rfDa4OFaXCmaolT6Sca1p6aG+t6dmk/JTxEUIm6anJBG8Ki0IwxUOG6ry9oOEVPPMAYxAf85
kFqV0uTbFGb7uk5FYUiN1M+R8vrc9biGAjTNyomX2ngvObJagOkTPqsAVxMgLZpf9YP4UB675cMs
7slXYjjjfRKMpkPqSIJPo7k1dkuDNWK+pvFWGuYpc0wLnaEtx94WbfLxmRDNZdB/gKwyP+KSuh/D
CRIqP3YZoo8Ro7BYublNAjd3Qg+qLrgwH3gxCMNiHF/ArBlUa773xD+xi6wnRtrT82Ha665B60+p
+eCvUHDee81/J32NodNhdvoSmUHJ1CkWzqLkXeQO9uAwlvlk2Q5FQ3ar5sKGeMCO/QuvNbVQ66RV
40LmSu3PdEL5lF6YL/JmBy/zn86dUdvo9taYHK6U1GqHp4yNcbcALmAjnrE6gOTxz0txsdy0wlpi
xxAO+ty+GdDMw/rVkD5bZxjSNV1NfWpqJJrAXv2R1emwy+onpi/FrBvZA2LvLp1TCK1NRLOwhdRP
fmWXIZyeOttyWTitTB/4QcYlIJPvoMpSG3siITmpEPksEo9WenwCo7Y8ungyuYE2MuNQaLET8ay2
QTJdOEscR2MQIv5PVZmoBi6uNfbOkp8FQteuO1gCvkRz2ehDDcX1ko0Y+sjC7iPwkphYvVHGWTE7
liptcaf1OeCBi/FXzB7T97nUlNRqWisRAbBjbQTjOzJk63PoZdo0hm0igBUz3orQiQuBHZTVD3Nl
sZV57wnDO0DGEsQnbT3pMj1Bqhw+mDfExJdN8PAWYnaYmSaXYLysBhZIwTazHK7Jq83RrcU/AHh0
qcEA6NJTP70vspaBdcNSD3z3rgVvPBFhrNIai00HJy/GwNxub20z+kNO1VOunxAZIjNqLmlEZ5r7
nPxcMAESxWwzYtv4dwzjx5TE/sUuj001Z7Ru0a9lu3aMUysY3YBufMlD11IaHekdaGdJeVk3rHBY
8/Q2MtncMcv90BKtsmUjKnlW4HJVFLxGxoxNaNIXIljedi9aRrBDE/r3vaeJylpwfnnHl51VE+jJ
MkTptc3MXIRYDWk6SOuEGnJISni3zYigGNckp0dwp6YQCqaYIfmLrkYUsTRjgawlHImAwXhCRiYh
IKoILEdl2wQZZwO5J2DcWHK2zS31MUwXeV/0nA0VcVv1VPD/jBicoFdR9MrnvD8x6DWdUUIGbSRM
BYeAS4SnbLyAMlabtrrB3CGdf18DZtyq1hi26ZFUtC7ZH+gtSZaryTq9XjsUNRQWBRMlg809a4yz
RMobEkqswcUfO2+S1vUm00BpN1PY4f4qt01izVwENl5uf1m9ZxFAoXnb8TGXsLdPL/2q96ZfaYsY
U18YAL45/OaZCxL+FZ7Y0Um2xcuCwUnzPXrqXTLxeqqRDYacDbg/9UQfYYLuQYSqivV3qVl28wEx
qzSphn+LSS+hI+Lq4flQowcNwri6u3pXrFek5oud8tN8D5+Zyadh1Xtxx7EKrapUWE2Y+aFfOWii
MmOQRBisscqvJZ5lN0WKiz+a62ykR1I1fy0SfebpGjoGYXgDeOnIjiA9JiWW1dw+wjDOwpAbh1Eg
o6YHtOcSF9puhH7k1L838OXBWOqnDRp1OgDCIz+ByEHUcOirK6Lg18AaTVG3iqiaxOVmBJb/vzFl
fynL1wdp5MlJncC57WtA0M/F0YRnYu8hvnRxj1S0ZoTXKSsOQRQa27TFF/JhWX1ExXsALOqDJj35
Ca0yuFPgFfwvUAPQXgMUZzWCf6nGlCcjKoHtnPbTMhMKg7CFqv+Do3Dc6CMP4tt2VZ7rarPvlqdP
F5JwX8+7IpY/aWeOQQOJqZ0+hkk0ZLVFoUHEujqCg2UVr3yShbCDztqRjgHeHt5Cv0+WGqD7AlvU
qAs7LHe6WcjhkYYwLjxyBeiNiS7p3y8w1QOG3pTFQb6Ksae6DjR54UjwxLxy1Kii+k0/kMNnO7qY
HDalbHUx1TV6KnQ53fKwZlnfeZCAqane7GmiWTeIdIValj+EfTaA+GhIT4tBwFVUFaHFdgo7iwIg
rkmQPxzecRt6j8eE+S6we9OMpShJg8XMp8M6JCqus2eJTIu0jEkd2wbcrcIX/y0tdt8Y1t6tE7z3
isvRmeUikWs/syOt7cNF914HxmgPFIq/ezXR+drlaTsIu0P1SIP+1hSLZ89qGvYloV+j5KJSjKzB
U0KWKGvREawMOs6X/2Z/n1nKy4rdLb4Ppcm2Hpr2GwcX1BnkI4ovN0iDbEQFPLI0V+mzRQfXyIJf
uUmBGs/ZIXhgdLsHwoT1VGVpg5iGJwq5nUbFhcbDykoLc3kxNG2FO1a9FKByLEPWer/KRt17+PCi
q7Ld09rYXsOD1bG7rJ/k5u5H7xKgENAtuBv5yGAQcPcu/f0YxWncejckIGv4tYl73vJUOzROCpb8
Hqehs2JEFNOiSBO2NCvWLlv13NDY5qIuh+xhJCYo/ufjdoiPTUXlyTTaXtbVKx4NeQCNuRASvmID
dYL+7Fxje7BQAqPM+AZ5C+DJwSNTd1dZGtlRhRGyC9bWuXDgmAwr8bwQbj0RrH030LNlMXY0Z6SB
QgvGMyt4Pp2Yprg3YeOKl6flJsDxJoGUpIPbRyV2A/sp20qxbFc1k0pbgE4siSYzmk3EydzH9Pph
fgs8AkBCnF0vxErzWeBNaq+4c9h0EQQsrUsjgNM9ZKjQAuBE5PN6b/7oYCwMOdxtSuAew/OkOzbA
5SQhYf2V9d0EL72in8TWst0n6UYhVTkHkg8re0GcVrHlnnTGfYU0ctzz2A9/vmtOLvNqbG7R4Kle
aBFeSeWz9tGF44ImT0dxHxohJIwYiG+zZmFp1AeLxC5ebqVLF+M1eOYRW6iKJXhVgN/TVGU7cRb7
vh3cFyq/kEn89nYfH4ECIGD795CqvlJKREffP/J6QzoWyTaa5hdx3E8glxp2Nos0TC/GJHAh2riV
pnpsjkfKBksJbIyVjBtuwIQIms4QiKAbua1HgqJcfBlTaW9yal0617N/xxO1OU6LluuvQrwKQHFa
EVmIBzdlwbQ2I+Im2zkeYfCShYOfFNXWe2rQCFBrKicxZ1h9/jDDPKsBK8pK3DOwsVozQg8HJC8y
ZrTQZhu+xknWDqjuZ2l3x116x5/znY6m9djg83QpL7cy/7IuCR4goKQp5GGn1maTzKps8e99xtCM
P1ki4qH+Oy4YMnMhBWi/aYLbGmR5tEkKyjdLs2+MGphmvgKbDStbuJp0jAQ+GpxdxsLosDi3v6Yx
FDTrIcsGyybws2xmenNw+wEOmQvQJ2UELx0XZmlakdYSWoTwK+iTCrq9D6wCba3Bex216Kgc7kdZ
6xKkbeE2F1lLG+gx0r/2jYmxq9T+Mv49oxZd5mxLc1fPpVmI55ujvCgc0nmW4EBg7MHCL3sW0UIw
bvq24oGxSPLm4vNwKJPVoxUtZzeP0IUMWuToaL1ogkITboNeekUoW93R/UYNe3pyUujp3sUOdpXW
X+w8JWX66xOhLeTqyWtzJjhS/KFFv0zVJ485X7Xzaz85eALpYj9gbCNmgzU9KywEY+aIjx5hYWk8
H+8NyeUilmXiNLxl6g70yd+UCOS/9oJi0pWeU7oPi6bUvq3GU37q+DkADDvylO2ia0OJ7CwTLs2V
MJTInbLdIWjcgW8ovsxMVnviBopAl64diGtFApZymaOvtJVpAdjhmJrioPwia/iLTpwq3qjznugO
opvM74mTEG5VdpsLCTMWWrhoPDUzom2C8TI+jX2hQHmlqwurUD/2mOIGIG1xwFNnDglN6neLPyPT
cSJWFNKnXXl1TNTxip1gRTlTw1EH3n83wIzMsrAMMBltXpjxISBQOB8i9bG4o9Bwnc0jctjPwav7
ls+d3e8lf6AKs+9WmQPhBoVv09iBqGMgGDyr0mU3PdvEjzD005o2MsJD8g4/qdvgN+NDqjXaLkkl
HxHNx4NCpWIzg72jrl5UAMDdLCA8EqfEn1LhI1oPsrdqmpL+PR7UwDYeIQWgsP67D3LPn4ZfhsaP
j5d+PAim9n5FOTfrlfU71qyOo4LnRDXEA+YEB+oWguQLMtEfn9mgJ/ZDmrrkcM7yRuVFtHLETnh0
6A1h1JeT+gZrz6rFjcUg+Rm6QZPlSdXtthy6VDUFZAGFqYBbDld/iigoIYNS4gsTJOP604l+5+/E
7HxwRchk9wvTP1tm6paElG2TlXhuOaco2V199ZpQTQbeitIMxonKA4LIqdr+0s2RivOIKVUx3pgX
I5dKxj6K6haa4rt2wC8Fx23ppp4326YRkDIHDxtrG/r5D7aDc/OjtrmQqbErG5gMMv++fEapIfxY
4yMEwe6hXa4CtJhNEDoMjV9szKoIyxJwfBWAldjNzWvqItJQgwrA9YljrdedW95ZZtLWeV3Sfk5w
QyQ/1ykeKSOeeW4csAdy34TmKZi9wigscNUmDh7MjO/uBk+r08ySXycIrzhrh8DrYyIlTwl5VUGT
8NAGb/JuLK0Hcmw3ciHmRJaK6sR+Pz97xihrCbBuLxJyYjPD0SCLelbrEYBKsQK0IpJkRhYiFDae
opswU8UKM8pS53ZQ1iFxoSK8t8IobvkAFACN634q0fja2Sq8qS4eEtCGcYHgVVvSZy99U65sh3oh
rx483WpCYER/iRgEbvZahnMLb3FizdzeL3VGeSJjk8ZlJ5LUO7k8+LBmIx3/I3ebnvSPWA60MIs3
3gMhsSYc8bT3ZsJnH8uMEVQ+EAER9QoGVeDmrW1+hlBeGmriIAj5t+GJ8/uhERIvWtShz4NxcQMj
Wm0efi31jj/MphHRPYW/sdZpEpOkm4LRlIPXeYViH5vhvPsEHRirydsag4xWYZVVsyDQgvTRhuDV
fpLlQX2m/+34Tj2oJ+D+Gtw6u/rmUZeDU/Au65+/bb8Gl3RTuuO1Qoi4UJdJFqVlNV8nrafJ2HiV
/fhMYXjMq0ti5MN/ulK/oPtX5HTN7pRLO/fO8IIOsyCO4Dfmo4+72Nb4aUDomxgiQsUiTqXbarck
y/B97tIKfGNSAJ6hZXjoNSbhZnyzzkc8gyVo9R3ggdtAIfokxV+kW3UphjDDx7bttxjmTZ54iWKO
hOirQfU2IibizqfeqM2ihw8eq2+Rgv0ay+PKnyzI0UjMu1U5uznozsPbLzbZE/c7yN813aTtUshg
RhT5bbAYvcuQcik8Jet3HX6xaCllgmT23OCnptHOB+GIeXyELWIGgwamolADO4qGgs3HJrpFu8I2
8qRJY/ZFgRIAjO88xLcc9qVX7OENg9rtqMq4pK2chvPiK56PSt2fQpAchJ0qD1qtOip8tdexyN4n
MtMq3xT6p+e8FupuQzIXF0M0uXdElzsy1dxgNec43oVTwjeynBkmPBarYSXD7J4/fweyDXs2w+Ia
faJkIS0XkTrXw0nqUv2SfIllD3TKOTMBim4QCNuGW4cU9XNmLhHziX+bkHCEJhqg2geDefYcK5V5
l+5ElcW053VujSL+kvFvQE2VLnrj9bQl+6uqrWgXmRS4enZ85OlyqpG7jMNTf9AzzKMW9dFFq4PH
l59jN2M6/mGtFlQdocatqiEJBtw5GTQmGXQpgSSko+O55CBYHkAAUw8LwoEjymOfJkyQjRD9pby1
//5R45MeIdsW1e0n/go1YimHvqHi45pNZO+dokH4BpJlz9/dqZZTk1m8YlIat2ky27OM+G0MFnyE
Ls9CaB0BgHYz1cQL5IDUvg/W2u1YlkIjHWha0YTi/m/QBXmQkIf0AJhhgZlohpwmlXNQBb2PvBnm
2yIQPLxVgqyWG5AT9DmYTbUBFRDWvg1+u8rZVLRzswtE6WvYSgUSHe8sAmTuuje5vdKXfSVrak3h
AXOw4vVYw+hkxCqy+F3Z3/N3B4A4BXG5T/eXOmHOm7NpXK2oz+dqGTd9/NbqAV//deb83d9lUHNz
xzIg15xlMUdZnEQ4HKMiIQXRYVByDv7OozrXkA7vNts3HEqqIOpfFeI9WyOgx3BXQhZM4rW2IbAN
3TouZNDNeuBgzXaMmzYavwFAsHvZxK0KJFoT4FoyHE4voiEpIZB8qcDLDnJeMr1toPVibr9p0DRb
ajk6s8Tih8U+U0nKPFaILvY0tbUQq0xZGoukZTbIIdvfMOmFkbph8G6+xLG2LFyxGn//TIyk3PZC
HGCTr2xF1LbICLh8CSsb8mNLZye/ABO+l3oqRLzgocTqXx9grf4utFFvAe55JnwbqzGgomrPPgdJ
IyGx5BCMQknoUK5XzXafjawXsqEfSTBGJS22pt0wazpIAPo00LWuadaHfxDc1pqEqjH/QVG7gxGm
175F1B0A7RJM2b6Lztk8QtDUYQ6CaRSRCqHgJCZkll3Cj4gDAGdEu4Mkwd4Nb4CKdtTVCKbCtlu6
joCRY/JSij7looYakd/bUAbikbETbMBvP/F4qL1DLtro9rH6ZhYGZsMz2Q3IGTMxCmUZhFVjIcvA
RB/02rxzeeqfmQGwMWjQ/VTJG8sUnXPQgJ0uHd1gJE4aH8JOX83+An+tYWcch03mF9M4T8VxAecu
+EzVMRv1bNUwvixNjfrQZsag5i4oKB3TN1VqBnzbiKz+yRfjQv5JFN6rCU402CLPIMcB3GkhzqZU
Mve0ckXdp55rAxjyOnehharTfKMHWMZh43DWmX3b74XstTJOl3b/xkGpmMLg+ZVGB+Ij3f+KUD3X
jReJ9WSn3zyNJ8kSxJQAXXRBFIaxCmMVlq9pIxAXNW8qPppgqP4tURtnrNHFsGmv/G095BZ4uXYe
ZPqgy58I0Nh32TjKh8Cm0rX7iZGZ7ErevvCCJ1uNj0PWV+u9UMkSGyLsh79gUGNZiVnbu1XIKNMo
j9yKz5bfOpKJ4PU/07FEyVytlp2dZbOwxvIwVoaEExyDjZcT+KyzPtIicd1C4oeVhiPtiCfpaYMw
+nrGx51HQNkvXDC2D+01rGZXVTdpz3WwXQKHxOlxfxLf9RTpJtRTacT2UU1suzSFiXRKvt8L1MVQ
bf4SbYIhUbb4Q5Kvgs0e1DRy5lR8jiwpnTv9K3XGA1/JIg96hqMNVklTruLYc7hUhAMTMYW2eZeS
EyvTVEnzZh4fTaanEKTkScDA0olMBon979NktRqkRXxGYBTymiRj7RVimkmygNc2xi6T36NuALhT
Fswi1WxZfjanYMrTFX0YKkOrN29PzRH72mii+rcnLEIPGMQAa2VJaNseSESWeDTuNGsJFMN0S/u1
WvfOi8wSzxgRt1Y8PxXOXDHC9Y2xlZ0l7zSD7AdpP7tS8V1gers5mlE72tKiMMfUS0lg7f7T4G+P
/GuYnv0g5RXE/6xW79xrlSW+oQeaqr806CAzB9HnAVSPFXKxscJqs1k5bZO2DSrPLRMYmHIuq+PB
b0vnNMPftT1XWMv73IrEW4Iv/DBhuywGVdOUX5lCi9w39I/c71FYcoW/mEv8gq8RDfN5WkWF6gyM
5nYMJNDEWsGc3iyWeZq/wSCXdLkmXKniEril2jn4pGGw3oldCyESfdCz/cDQlAP+Ki9OQ8XqD1xI
1mcs7PNeC67/InQNIv0Dv9nJ/bxAA+8vfXaInawKdREkKf63Ybu4tCT02nMp3W9edZXFKG5JYd0N
lInVo890Ir5Hd49ruyjb9NcfTAzNN6xAeZEInlQfUaVG8C/KEvr90osf5RuT9filverlOXE+BoEF
cZJrUyPDwuCF1EqelIdhVG8rlFLk/EY6KaaYBZ1ab/cOhh5Su0ZqtpRYiU+OB7ZtCph0sqgLXvwv
pkiM5+oGuT0qmIbba/s/4CR2JEpeVvu4+HLy3ga5WW5HdvVPRNBKhHtCnH2ku79wl3uEEWsdbIuA
KQBGsUL0epxoU3rT76fYHJ7saganNf9Jrno/QZd204lwn4GSXX7gzql+yoobNZaXMqAU3EIqNdy1
68Aun/6Khuph0oX5l9iFwI06DXBbVLv3e8pMcD9OlQJon3fbBXxZds9lL74uN1Lns2iRh3gj/BcI
VaWjZChGF5pZLUbcZWb4HZ3ejOFs0QMq9lTH4KoGyJZ7+26rAhNsbO1ARUt1sYBmoB+WkD0XlDQj
o4Bw8Lx1vuqj7zaXjQk1j9nzNAleGfgc36bLnyy/yxcmFJy2cWsVrJHAQtTAJyQ4xk2DTx8U4AgD
F6ZR51xdA5h0mxeWyNu/ygqkqMEgxhUJ+y3lfDmwFHMmBnWzy3wgID2Lj6KYEXqufQwhP5wZXFQh
qqAhQwrsiW6Kv44FQcfv696tGFR2s+Vap7OKg+u1zxeJSecI5Jnspop9AWjrW7Nvi3N3ndQ1Io9b
ADUsuiKAjeo0xA8CfmqZCZIz0lJWc+ccfQPDBhB/7twoBglOYWgDWCFqSXCYPqKGzl0qFeA+wey3
140huv0qTfqKIzmE0d/c23WBOq1xAxkUiJ7zEaXntur0Wh6X0L846INHjEAJpS4NfQE2QBn0qj8F
RYfKDziG52Xi2FGIONgN44u5QemAZ5TW3sm/X5xqkQhzuHXYS3HROmS22yuQY/DfDsZ4nGpvd8V/
8iCZJ39aFWmhNBc+TVaHYIk7FimZIcFofG5CuUq0JmzqVcftOXwOtp+xWotxCRv93kENCVSahUbd
stErqam5IDd3EFSkvlfq9D6huDtOkKJu+dVQmPKSz/kjSInEyP1MRDYosCxqbYOh5EaKO/O7/3pc
4KnrG6ymMFFrlkNnilVnyddHjGWHoRtx9fsjBbUTc79wTw8vbFpfrO4jOjPESeEJezn3KZtXcDtM
F6uJ43KCDq2On3vshEO7WvmajJbCcFZa/LM8LEVlSFMk28TzhWSQNwxDrFSBeCTiVsZq5CVd/Nd9
Lr1QOx008pqnkIIGTp1k5M7aXdggC2D1WdA73iyjw7l74u7a87Ze79lk3k3gMEaKdO0VtAZwar0L
Hm790fQC3VMbLjFJX+tAxDtIjT3Rzp2VAnU6ZDc0WX7reN/58W00+CNF+nVwulomDQBad3kgfcS5
MFYwacjRePQgJ032rnxLgU+43uebVlVjhbHVrhH+/7Ai3ntouImov0iB5+iKYKk7N4ApHB1YGnqc
vPPoshHj0lq+VbOEVlly1/1mM75/Ifrx4/xqz4+MFTC2a/fKIiJYNMeje/IU1FBosh9xCz1hUbOp
IjZ45YIcRCdKL1jfR/dRNdTvrkJibhwpHZrJCoL8cxfDf/3VHwamWewmywAaeY+n0FPp1WaH7o/4
rxp4U3GqwvRjCeFYVKy5MFr5Z/cOj3zNaUkEPc1TdOgKShEjyxvxv2aJKlOziawgcS7ugZEWntQA
GCPeBsrm8lkxr9MhyiQ76e+oqX8YdoaOb4ACxawRhMHQaK1Ox6qcTr4rgr/hTY+tuWf/L06BNu7g
c/HmsLTvYi4At6GP8D7ZFl26B722wyqyHJEfwDcNXdWJuJ1Wup3ZfppoEjL5kKQD2rfmsedN2b2A
s1jEbgz7xotlurSkmJBDdb/ueHQOgQ2c/rGo0nBi04EsxOFiGfKerSpwt4/bVtI2UVLj3xsMwq23
GADai1cBQvwr2VWP07IPQI1NUnoBdAh+JJ/d9KHSyBUzrteelnVvC/CfVlQ5srHoE2iEAhTSDgLD
DCbjlI6rZ4Et1DlDZSlOg3xmc1fTHaSSsAWfmFoIYBT9eIqGJX9Jtl/qCD1MKm+JHqH3TjwYYvjl
G61bjeNIMOpjFl9btZjXIUHtdhmqavJTw1Algw3LLI/S2r8zBkETVuwDRBCF70Vmbk7EbJVZSjSe
JQxUVRnupoBmrZ5VeV3acZ51OAE7sRYsq+20kN3Dq/mbGuehilPONAu5GtvKshXSnG1W5oGFX3pK
O9yvWI0ddxS57ylrfQ84DO45UFnY0Bu7Efu3W7bU4RYcdaceunjM4Lzikir/LyRIMl0TVnzPSHp+
qk9cMZQWUMrgRg0unQZfF1UNhFCm+4VQFI5w18fKDwEtlv39LpZXbeWMMlROYFhLT/yw6jig8rhg
8s+N8yjO+sx0A44Eq9/DexM89kGn0zBmW+qPKw/ZK3Ew3BNZvIoFIm28UIwiJAoVchIQ8U1Vzg6g
iKLE+UavkG4EW+RZrfy+2DqfBOf7d68aVY+vwxznrS4jLjZhJEUV+SbQzqVGkxit78MY8EHXh6hY
Z1TLZ0pDBS7eWFoHagxjImcn8eR4jcETT/yFbcG308GvJHuezPTtqq1XjPYgfn53gqe0EFIOKdll
11PpkMQh7RHjoOpgTPxUnLiWoWPQH2pO9q554D2PmBgBQUFQdAI2snTbuZxewnBlJa7wBLxcJo76
ZjcJiNJmgM4+6T/4yuj2MDPHfT6q3x3qOowwFHfaj6ZlUuItoP0z8Sl22BkY5kjjVxhY2jY9583C
n94JFd6e1MoK+U/guAO8iTnROibVJTuRVgKMt5D7J7wHfRep6xYg6rQXx0+RexhPUeuuVqEN8ckW
WsrEYT3JcwxOY4YKP5YulucBdXxB52SodX8V8l5sh5AlThKwohcwBSczqOu81YLoLgcOORTM56MU
rhoYSgZWmTVmZjB6NJA3Uk1x39ixPKHX9utzl/XHWx021aVp4Z0SAn4+W11+3t2W61l2X2TeLLQg
fbZRIRRl5rCR0cVdHFqj6cXugHwvezXsbjo4Y5ZuTRq5Gf8HX0Z0QePSccRHDC+chaDgXBfBm57u
wv/vp+FYiOCVaVi8d0FeBWH9gqvKNmT4MMl/OpTMLBYCg7uZJCZ7j+vGeEhSRjv28fmTMJIesm3d
Vih4tz32RBa6R72CO/pHFRZBf0xWuqyPvzX/M64r3ntRS9QDf/ovg0jdXpP/oqmRZos/0rp9yoMB
jT1bRmWfJMET2C/KrIPEPQTlGW/4vn0Z89aThy+Xf76mAdbkZ56Kw5s6qOxqte1S4VZOHHEcxzG+
HJefCdZXyzgrBImaR073Tij8868qxYSmcNMTxzDip12H7am3S4USEgbAsxSaerjAu/gnYUJxOAwh
PFWHecnuRvPvFSBTjM8omA9ENcK/xB3CRPc1Yz08evCqP9AvJMA6Ix36frdWvGWqvL1hxfqNSoJC
g2BSudum0k8Keg7NIuIrP4x58hXngHorC5GpE2GdBP68zkFgRhrZ6W5OGw8ES76s6Z10AxVHngTq
jiDR+LwB2XY9iP0ngdZQV9HkyQcZ/Pyhyhjt1RhEOK51HIgLCSSE2XGT8thlJsZA9uFx1Dlvwwzz
l7V5UUkssg5bkaPr+loyF040e6IQ/9geQWcyHMTx16FSqU76mXGPwwFYdqF6mf2+773cYMJCE2k+
qrDI4Wh8TxCKE0uHB7YmOhwG/puU9JI7UfVx0gC4ORAEZ+3otf9m6olfyDLqR5ogXMSgSz8lveJ5
QpbtGmIaWvrFgqgMXVGjLrRxN9Dy3kYKaF6YVdbH1cEjWHea42Pm3lkUN6I5Vfn5zE55IiOn3ebx
A0EZwlG90wtxq+eJPt3ntpytPyVMrXpJiCXt3g7KBlfMouRfPQi032B0sTJNeznypAhL7tlNxrre
r4Ddk0bSd4istVMvf0wgPjtOkYtuUFgcPoJ4P+YIAWFfixWdm32KLgIQNq53Xja4BHlIxlCvhH7H
A6/Hf09fU02zH9hPEvveituAyknM+dlKsyWyAUNJ3qgo/aSSM40KcVOtDu2VpJFit3JMnindNd4A
JzDIKkbVhfuDsYg3+8p92VMhM8Vz8BrkW/cMg82EyXxBeGIyUxaK0hk2TAiUsMlFX3GsIRJE87H1
p7xOltKHIBLYb0TnzBjKU7FeOpFaHVFc9Cfoj8nB2bQm8pFdRAWsBzlIZ/H7HBSupW40BPvw01f4
LCPSKff2gR7JLZb8T2OJdSnbuSzrl8v37yrnKwBbGe+7yz1URe9F4xL7CjH88Mperl38ZiqrO0kU
MXwqE9NFPwaNTU5SVP4iF+J1RWZMIpcm/rlLhu0QFBy4/yHtHFC+QdNYh37+DzXNKaMe9Uor/auy
BXu/WNsPMhXxX27bE+BcgJ1sEK4kWpo59kUz1WgF+5mRriVYVYQHnzas3ORaHFVc0cgpqRbnkWi0
5kOda968C8GmjAvBHHSlP/jEUxqPLMBLcNBs8iMoi205TkAJwNQTMFK8HlRNuy9HRmnrJ6OzDZv0
RkJFLzQOR3tgzTOHm7Endx98+7SLQeXWjBpkC8rzmk/w5il6JH3wokt5Qwi7hBMH3XMJxiXCPAmR
hxky5jP7Q2X0cXvdN2GGCxnYlTk+MB2d042mrmuWjLLYdYMBfE8svLxMcmDQ6uJnKyMVCo10vVZd
cshnYRkCMkY7ErQ3ZMT5s8fnVZRZGZ4EqJq7c0uT1SztBqC3c1TMyRKv7tRebCRWnQHI+pSeZHge
5ltSwLUzyb5JigT1JaYE2rT9LlT8P8X8oaB72i2MYZier6X21iCU0+9dju8GnJxyB2fcRY7qVa/D
zeQpfkrcaVFdGZeSLIuS8Q56GkyBXomGhPWIWfdLG9Xk4exHTz/i4b04AvJWz6qLH9oIZTpPA+8I
lBvEVhMXV/KcWfMOaO2MutYwcdP2tkEfKldMHXFX7+9m3J4H3e+cPXIDoFCycd9ju7ogrfSGRE/e
3VYfc7cMaQ/2YJ/D+RjkZ8a+X1uPvsKibisgLcI7sQyZEH9i3t4o0Oizv3Nf3DHTKdz/3bLkbUIj
M+SLdR+tHJS8KqVE2AwpCSdb8qUppTaSttdeCcaXiJtYiuR35aCYYGLB5eL33KAfRdKjfuo6ByKc
VukNFPu4RSz0gnNDTv8OHhQae1yE4atjFdulHx3L1qtKT1PCIndYtfiLzBUQAodQZM4mNgTSi64p
8eiOcEXoV4YYIfHd2SucgR8FORClNwMHvjwhUxzPaXDoME3C7Igg8U3G7IjLqaNDLoUT15rj44nu
okanEX6kaoHD5KCCxl2cKQhVxZAFgEEQ9BrnnTNZSuMR9+M71yV42kbjtAApiAyjhatEI3PWmsdN
bf9ecQc6QRsgyCG9ymGoA09b7s2UVD+dfS0uluSPXFckh4Dl9KngNdSsuokvwykQWNcVvy+aQDIl
SBPXV8ZK+6UwOB3u/QGU4Q9Pa0KX4B7M+Y0qIKrFdsuaEltehZ1vZhbv9tulGat8mKVikP5Z38Bk
qIBBPnONPvlBfqmA6tk9IzD7WD6j2fxUXiQx6j4XBlY318FXTkanf7C87t2rbC1S
`pragma protect end_protected

