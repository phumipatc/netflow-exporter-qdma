`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
g7xG0LGZvPzJ2/FqokR00Po0LNGUsZ383BH4OwZ9Vn4BRwkXuHJvuOU7ydAah9jUV8Q0YevEqwod
9VVaY3FSP4+QqDZOKjfm19gA1MZ8Rr2kTYqukzNk+F3c7HM6V0l4GY+o1v0oGQ8LGcTao8j5LCL4
g468pg7aw2qCllKTG6XpJz49UzxzcfN7pxKYPP0oFKT2+yF2t4iNr18cY6NOlZf5Id40zgMXQZ8/
Ozyk3DT1F59gt7gZTIgZ3nnHZUfMXbswKo/mC5nk5WbwN7nYCSZhbiWPauOZkLqaXvH1iAW/7qe+
rtD2+DOdt0rGa/kmdPuQ9Q9NrQWLqIEWp5Klpg==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
w4WQhDKxchY/uWiMNzsQbOLzC1WINSIMXasQ0ChkRwpgUbJAWgMEJJcBS2XHUT5Z9cmBYHn7H/2z
FQGFC8MD5g7yrjD3K7tiFCv3NLY/fAARFXD8hjwVzwVwu8ymCqDu+gVp+oeihdnU6ri3aK4GIwt0
/cfrQyuZyX1V+R+SUXESkhcez+ahiDfvR+4LMKYgiVYPmJ3n4nVdauKr93ioIuLOsUPIg1jKx1G4
E56awHyfzPHZB0tgE5R8CE07iQ3IcXE05dtjBEro4M4xsoUEuc0TQL7Ah/v73yR6PbGXaB1WWE6b
bUC6ul03ySHTGOncJWQZFfssMZdrgGKyc10eMgAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
RD8DD46SHNheO6vLlkajr5t6TIwtTsX0sVCGr4oGhq0OqCYSVva+v6cdNiNPzwEMz1Oljvz+wDVB
+p0WJ4UdRw==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
iERytDF35AeqznwvvHoEWYuCAEJtJ+VMhrqKBQcZadhi1QqKY8AhRw4zm8rAYM8qvd0rF/WKiqfO
hVDdf5lpGvWqafl4704Bh+xtsdahIOVxPSkkRkswKU56+q0o5ki9kduN3V4QRgqZOgwZ+le+fUg1
K1XsWx5XMrTSyvR+4bRW70ztbaIjk6nWmfvqiB3apElyJz5HzTMiTFlwCjtdKKrTJCpxQcZBhW/D
QcuIWMTu5QxO69kPIWu1PWY/yMZnGbLyJT/MnR5qEVjLvpfum++iRJ9Ha9MPfVxSUdwBdoUS2YY7
IjUgbJxQR6dUeOTEbiOZzw3T50UyQmP0di+33w==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jO/L3GDwQ4WJ0r4aixVj32fwvHidq5UdHwOUu9SrUzDZFM9Oe7EJnme9//gnGQSZ2KT7I0vSq7PS
K/s556TzGPVgtbtDUWNzQwykhMaCdLzC95VTxf5rEvctaszeb8nrtMi6IqxdaiqBhQ5BDwwf+x0g
IFSBq14WCJs/VGr4akjv0zkw3dpueBTYhWJYxTqOy93E9TekWlhlw1tnQ8dRfEv6NRRFHLbd8HPG
0EbfTtwaDUJXGIZ5l2sGOTDIlCXypF2CClkSF0IcfF8XwvwtaYkZgoPVFuRAnyFqATm257v+U8Hg
WgnhdiCp+ZmQD6NnPl9wEwVYQ4J2OKQI6GsKKA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
UUEhePAa4Q6+Rk5SZiWyQQlldcb7OAVYO/FX8Cg8F2CC73P/hlYHXG5IDqgH9ESiQ0fM3dPZYpcj
BrdXUkNAh8VRpYLvLAGaC1PfAQXH7e0dbNvHJtMro9h3mLJ7Rci8gwUguApMFGNW6xMhAc4GMvYt
MML4QAM5LrjHfW/h+a8=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
UNxEfhH8aqEpjfLuIlv9QWGchJeNYR6fDB+y2tujUn9br2l7XWR750q9Ldn0TX434WwvA2ScBJUQ
whhP9hg0DOHF8oAMZd2O/yzW0daD9iiJVu32O7Iyjn/OdGpynTIyxLSiXaBhhAmWDFbi9pGrZ3LB
1WyhAm1oJsiRmrOHl/B7OhA1QlS5pMuzWdTH8fcoQhuCxPhDzXSFn93lqifUjSxlUJK8kBXxc1hT
WdG5KuP/4eRzf4rT9tmvEJL4guWM24MuGNSPDhDEJMQL18D/NpGltD42eJHRs9zpds+s3XFaSdYq
JoqsqxvphdXrkDgrhllfrtszF9VAAhX6+S26Ww==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kKn3LLNUId4ktj0iMPClrV6iBbl5gU/oQ+/j2/olWSqxygmkeCrFqbCncMb9jgisGpAwjNmcvV8b
tAeB2MPUBLSAoGP65iLrxrctP7+x/2DImLivvteHFBIivuN5MfKQLYKY5TAcSHSM83O2cLaqpxgG
HoWfhBOvs+A3ll2ulQZJXqkjREhw+YGia9NAJqJgScOV5/9+M2xP/Ixonj8xOWmeCh+NIu38/i3L
WCp8uYDCJG6Dp4rZxkC4sQUzzJrOoSY46JnZhTjWZigdMvmg8CKvlOwieSM6+5CV+rg8PEL77aLY
OY7idPIsvqJainV3/1lRsg/lN/u3i4EiRUVTeQ==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GfTyPTZgi8ZV28IJLrobeb6JcmGmtlPZEZmCR+UZeY8deQv9fFzrY3gjuNjQ6th+mHQUKTFoJj7M
iAOyR1TfQrZkwb/EkqmeBunuKRl+WP4heEDWoKmH+jmS3bGOYlWW8ERzNMUUHvfxOQBFov4w4kNQ
/vzjOGSSMG3dIi4j4MY=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ii+1ErqQq4ufgvawV3LWeSpdEhJ21hN0xMHYF1OmVZPV7yzMQ+dw5Nt4+I7wlfMLuQEbMxiQHikX
csm0FwfjM7p0Upzo91qSzo1yr1peoQBYUIAm8a2U1a52d8KHbofPGpMaVFPIkObXCtutTo0OUWa8
1jSbzPkHsJAnFs17nPPTlrduZg40YdDpZFigXPxyNcCiGI1gCiANNk75uUNdg47sE+5DyrcSaMhj
a3Uv8ci8kOjG+V783TYigRr5cK8S4Dc8M34eO35ZG7VXVN2TOGRHXTbmAu/OFKflXYROv4pI1jjY
KdxlESp55Qrz+WEOhTxupunZKOM7EA+4rmMXgQ==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`pragma protect data_block
tAMEe2L6Ex6O27+qmA516YuWuWbnUtZMX7I4VQf85sVhaIl63PlrqIitVOxnFhGQ+d2Y/TQq6UaD
kmiw/f5JSXmKRGkv7y6CYFuEx50KQQjoJiCZnw8rNR+/7CvnV+wS4WsntG5HVOlH0m5WS8vRzKDL
83+I203UzNPzmmz2jPP6CZU378RYV9zRl4yD8JmpK5W9PylpAE5uJIw2JRSuI5MOs7TxMOAc4h97
LhFogJQ+CuMkKS6GBIAIcHeOWs4KE+Z3ChDKeW/eHhidNFu+7qLKhwmLtkXRJShQm/+jiXHiRgXw
XiXlsCcCR6hsl6geDeU+I6dvgyEmt3Q0W+jRC5cFhHUvHwf6fwwxITiz9qoOPxzfjzv2Retcd3we
ikM96NVhibAsF93NsjYOSM3e86FutaWjRQ49hIMMOxjkgBK2PwE9Vwv4FZRBJ5knEpd8ZTzgyNWq
oB2PgGKR2d9kesFYC8ii8PzGGGDsd5t2E/lTECCT/t09Y+IhHWo6zE8Hezyc6rAfoIjL9eDbQR8w
c8Zx7+5pWqxLNTyOVYKGdOKjkUM2ytBx2OL7v2k07d/+C05lWVj/TZfNqImivkOQSXiInz5JXBOR
Ke0b4uV7wIJd3d4vigI2buvpz8jayGCLBzbDo6Xupel+2HSZL4ic6LuTBVvdwhdLKCbX2c9V2/tT
iOzIcbXxp1aOec18lQgEsVbRHbpSSFaCcdevpi8zwxY1VEzbpYaqupe3PhauianapiuftdkydNpX
qllAKyUHLejtL/wdZKt5PI9VRJcVIZqFEfPBePdYC9WPUa6tnqPaAEQ3xHpT3NvrBkkND75OM33S
Mehbdtc7NGOBu9geSiGp0a+ZsrFgczFP+7oshqPLiEJWVAICNh7K8wYAua50DuY4qu/kH5kh6WCY
P2OBqZwu3w+2g/2wSRIfGsFuXiN0rIf4u8P1aZQA0k5cHDiv613yXdflm82Gm5mFLZ0CyxhKNi43
nJAwsfeiUgGawMwKTbEXYWAyBdcjS7dNlbyA0B9ofnCiGqYbl9wUzGXxn3dSQFRkRq/7P+sXC/QO
OnfzarkfQodOVdKW3gr/QjfPouN7PxFbX4fvw+Xc1Yr813OecR4QvjbfHuGk3/QdO/0ZvxDLRclz
Ei5tOwT+SC3yJ9DX3xynLdF35lrjTkrMw1LXxt6+hHYhuUikTTC96YjqO0dG5xAF2lJyvzC5WQya
c1TwreI2tU8TEwW4eBi7hZBbQ3T0vxFyFOy4WXJ3PPKWmz/PuBuWar4YYMn+CW9D+rHCf6jofZmp
GEw1ci4BJT5y7sgoCAChjep6lOFVVGZV494TkfY0jTVAevOGxgzsKWnEDx8RmTT1vpP23C0xBkEE
MEkNkVi4n/8LOz0cBPE7+v0a9L9VEgQaBtjOgPYJcRA5o5g7YuQ25hj0iNamwnUsKw+kWyZU8XWk
1odrKtF9ngZikmFlFrlC7j2Q8gJXdu/ce9uDdUYbuQ2Jettj71XZvRUmtw+raxZRY7TS0DwAyDaV
d4NfPTrQif6U1zHnLm1I03xE4Ul0raMyFfHsR6eEulurf/EYKhj89XeAabWlwACMbLZrjXNanVsj
umBa6OE+KEItgXJ66vYE6FJpLtQw0xC0zztyF3Y5Tc2fjDmgzLkBul15gGZjMVwNVGzeVj8hc/FR
/5929qYCAwSFGne6/ewwrWwJa+Jzf5j9TKoHKf0vCXfl7iUFYbLUz3Lu1WcUK4FZA0YJls9JY/yr
qjYLCZvjigPwVZViQi3iFWi/kNy4VwXyzk8cmGyqG/fjLSp7uGXmweE9fodraaLqwDB/OaH6QwbY
Ykd013tb4tgrRMfOMG6dJjVTFHzgMzmmHTModG2vEnwDtG7hgdbNPDYg2FmhAenGexWGnhzwYERb
zJjUD5TgnJfQafaO4Mu5shLiajq86wwzaJJtLWaqEQ6EgJx6XSiypE1JmexqeiheMPllAABRmypN
zfbXDrWmDmLiJsMse27UG2eIALx1szGgkhiptSmZr8OCGgL9xvC399ITUecWQYDZ9vgBElwlSMEf
yRHd5wBHCfWC2AmH9SZOZhLnEHMTD8bueLQzkkgM+9TMPEvPdWchwqSEwLwqUyJ5PVfQP9bc85cs
Z1gBzOWMuJ+lOc4hICqsVxlh2FtyzENP9TPx4Mni6x3u/miyOvmdHwZX3/CeOU4EBtkVStwiSGqC
qRreEHDDq4hxbDTXgBR+2qFnZl4TGQHTXAS8AB7feK8bZ5DrfFlsT8tb0GaKHtgsEngUnLJDt+zo
QqyTabp5ejZ3/mXQ5iH2UF7o69QgywvPrzM0meLnaOlcvLL3aXsHBEN+OrXrfXe6TFbWOmdq1hW7
37eLLh6hRtWoSPAd/ajjkaI+mgSLNxIS8KCzJgznNxpQQIaj98AbMUGkHjWwX4iTRdyiZlrpBV1q
qK8tdNl2nYspE+ufjVZkjuOyZeTjZ503pgReByOFdWmln+OuGLznEcoG/pgPdlk8LRlP3ubVSjml
KcUdQVHOqAVaWQOPZ578ul7DxrO3T64a+CCY8+tcLy3V/NLinC7BtoiCexvdEAdc8xDeK+mSXTkh
SaUxMBVuxjJk4HjMNZ4NWz914MncwDdieYTFSp8nxhxS7zghPk/96MucR+SwK/RtQHRBq5WU4FZP
+SMLeUrR0UTCaEfrnVfGZ7TAOsZseOHr2QNsujzvLH48GpDIzpAcTY3yNZ8NRx6vb2QVC77kuo1R
cCxPtfxxxah3q8nv8KNvTrXryN6tN2Al49GAHP1Rk/pM7osmJ2nIHsKPEVLETdF2069V1Bsh9bVc
nMxX3yWH7/f9kAZI5M3bqqybzK5uMb++gGVedDi7q3xyadhKXK9/tDVU3FG+ou9TPxF63fT3DqvR
VM+PbG756JfQA57Pzf5kVKt/dGitNB263ko6hqhr4qcsio1TFFiyxTBFs10L9A7brQyWMbjnA41q
6xQx/3p7s3OmoMqTwI6kgIJ2iGcYUqVkN89RWqK0mIJiASJfvy9f4ezk9p5EL96a1m+d21UWdmvG
Ak5ZzYDCr8zww2TERHe6PM7VYS4FSb4kRm0GTTm288S0YVyqYJS8dVDQOk8+JKH9zx25Rm7RbHIS
qHxy2TyxnlAm37DZs8yfLnOd7m1Wo2tKsNG5/UnZePudfxXEQJ5EOZT5Dc5BkNFcqDlUuTtAEyGX
s6P2P7SWxTN+hbPIuMEkgZzUDXGKQyYjbqTup/qQvD84ggjhsd3xEU6wPCFCVg/347/jZ4yeDq0W
7ghumKjqm3kLDzFp+9oeg5d9AxNyTHt7l0vf+WWAdHLxKoSBMB5CMxLpodStJ7OqzyVtgv+ikQ99
xJ1EHeKAH0eoF1GhB+mcTFuEH9I32K5XjRIuh7r6R4LDPXizWyO3JeJO5oNuIV/0J/2x6ywkEJld
27K/dqdEaWR7d6v7O9XgtxgKXe8wPEiVuycm+1op1chAdHA3XhowiyHOfjiclTeC0Own99T95P65
VmTjUSwhV31wnWub0xBgj1JW2ZeARiu9Ku7vOdtacXPngbgrJaCryzz87m6r9W6boiS2Ld45ci2x
JuB/0DwJbjzPo6jAOWemVUh0cHh+P0k9KF3Tdg/sul9KIrXXpb/nSuB6ug5YSY4aB8M7S+o8UbTf
68+keVPxSjKEKr/cgP1Jt8EGz/m4/aUf16z8rwjv9ilG3D0rJdCEJw25AC6IAA6lR2ZYK26FF+Vz
miEjX/qdWQkCg2Eo31DMd4dPDIum7k0FHsxt7ZvbWAwZ+4TxmA8Nfg2/sTzPoRqDOqUq29ymzZre
9utJ3UBJZA24/wgRuUXa/I8WwQ+ooR9MJxzD8UEF3Ca3GdQmBLx9KomY/rZZ1FqsYFvlPmeWfDTc
kt1eP1CqOsskgKY/j6rPmxamEzMbmJG387T1AO0Ka5WIKN4NflXq/8LvDvPJlihOJVq1FTs/lrUL
7oTq7yVNpNa6luX/QujajR7rgs5kD72bm0utpI/yTq2IpMW4bh3w+ZNMaB4iCHk4cKhXeCFL7WwJ
cGM1MqV6bB4H8nlrNBDOzSKKYQSSkzoJob/qjOorWijMk0aNnN7Kyg6I73M6/ubv/zN1T3u3uhm/
Uw+2DRXmGVu5PAm4It6el3nyBn4JUr4GChYxbko33W544aCsvCcwCssGHksXcFnF1s0chP6C1re4
fI3h/R71hp6luDeUI7zEUj7QWirlG51bel9QrpX0Nziu
`pragma protect end_protected

