`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Xe7uKBsB3poRUxaRjf1yX9Z1mZKw4i6zl9S0AzmUN5yQAQOuZ00QLR6DNjQS+9hjoi3BACdeUnU0
wD9SHPRzaCNHZoQs1I1QR/KVk5tNlDXQWS1WESL7FBozBsIhiyes9l6ylb+Lh1sNWJqycvVhC4AB
E1JwrIwhM67wg3be4B3NefmCwWN3MvPEFeyKV3IwEbiEFcOvYxggSPmYVIUjy3Rz5uvgf03uy4yF
HxAWpW6y9x07yIRgnLd8YqTNEZL6mAnatCrQfZisAeaWSlVxAIRcCuj8CPSAOGGzojnGdGQy/Dx2
K96DleY22ZoQSYm2CNN4rBhi8E0kgls6xPo62g==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
ya4GbFxttcGkypBYCo9Klg62yLOOoGDkXIhaina13UOYpbs5W6n4bFWTl1UiPt8QxTA7lc8/6twA
eVvvJqMpP/GLjt+myOR2zW29mapDdXkBqRlIsEzl/9FT0wAFYFv0PC3iEi/XhHEqTOXb70Zo1TRu
H4V2rEwFISr/6Qtes2l/tTkPwUfpwYkxXYHCR4oEqs3ZAfRh4tSylBFgpEkw4Zf+8s5u1gIshFt9
2zjp8TYl6f1oKXmfxLlSIXqAyCWRofGSzRey6hupE6SUsMSShRvJgvJhJDCPq5OEkRnAc+jMn9fk
/QdYkvc4ZINuHmHvGzVWR08f6IKLRxAJKc8H+gAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
eziwV5kZ7ar8Eu/E7/BZZ4r4OdQxbAdHM8hsF6Eo5blkMgyP5f++OmKjreLDOaw5n2ziNdajtm+k
zqm5fHtP8Q==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XIGksaeTahyZn2Nqh8zhQASLzASYa9Ju5Fm7jDq3RC3aU4O90X5t3xcfxqB3nGaF0DlD5lGL51vX
BaobVxjyHJq8YPnzh3M/O+eME548OpGadaer+SkZvljOAOJLKtP4aGHt+nl2/3XkzWu/to8i8mBM
BHdBQ/DF1aEJZNvtrm7EJKZiN7IBnnAqz92G0ShdKEe8qedAhXCYy9cfq/9RYEZbnxxxADBKFI92
LoVi3XzRXVMlurW7nmTl8Cd2pxGVykoT2fRJK5hIohaqzPlJmG7gS6aX3yF+1B8nuIsIJiSDEo6g
0iFZhqqn+Dg/Hm82sdLV3I0KqyQPHjbpCjQzYg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rjGYYfld7iC2BQt7cwJA3zM//2xACdG72TSuOICnJMeG6KOSul19QgkVmoJtpTSzPrH+WtW+ItXu
ZQVMIydm24ZFOM1ygvUThf3tkfCN4QaMk1LaOBNDh3Ip6YvAO7/lwDO7zQRBBQ43/AZM/zK2s7yL
qqn/MsUqibF/q9DJVojwNZ9u9+p7PFK87bjQWir4Np+7Lb6mqeXWhZoo7KnKI3GKQPgp6T5eUqyK
94atnBH+LW/lhAQyYfNkKgBQZj4d1vMtMr5+wmgPBFkO4Xblci6xcm/ezX6y6z8FTwOxJfe3bIaL
ilI7OJaSOoa0Gpz80OqSNg/2Y3Ud4cLZ+jY60Q==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
bKdZdM5tXj121O4wM98aBGBpW14z9mmK87JgBMLiJccdVhYCfP7tP/J34YHMCXGdcs3OA2ddJ+XS
WfLvHnCjGYH7NZY2ZPGd+tlI9x7VnO4mKomfM7ev/IZ9ByLIE5Q4gDZgHdb7x+3EUsRJv6/aBobz
shnotVvnUewcN9yFKcg=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WBPlvz1FcSEKkSo5mNnW9KNmYgVkgR8AMCoredGOy0+xAa991kSlxecl6YTK4LRSOdZRNh78JZdC
Xx1KMWjt/8qQLXhRdWv+fCAbhdI0PjV3U0gIdvzlAhOvj0XWYCdnE/jUUZS+DUKNFTnxrrajvkTF
TOxvtP5slYEYM0t7WSB7kmBzKUlcdR9BQXt0CTt1lM+Y6nUbLVymbpcnKiuyqdls7TK/MNgCLRpe
fKiaecdou4Aaio85n+XRIL6i6VX25vMMByOfsPupKpy01cAgqfSmbx9iS3xnvc7KHPEsHoq4wBdF
7ySDR0eU967qKqpj6SJpJPfmPsbzl7BdtA9pqg==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
cGiXZOI7p39XYpKFCljs8HPmqRe0ulitzgAFnYVXNq56+BciOj3jJ57GIRHT4duDaVSdTksaAkFW
DPtzKZDpKQMfJAO+d8JuOms+TDGj3c7hFqTCKWtWWYobJfbTB9YMgZLNtU02Rn0R+ZZ2Iodt3glQ
0dnKy+hlrAfvp5gtiCyQ83qQXKG3NOlE3cVr9W4PTy+bgz4Li1l8lFdXw3/J3WIy00WHNcFJrqm2
GBHVsOI55bQuhU/e5OovR/+KvcvRsQ4cqLaXgseIjFg/lXnlq5Xz5MN2nnRHbR4KHyEHMFEOkfAV
3Uo9jS1NQGuTBkwdwUet9/kjdhMtvrG3nqbKbQ==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
HsYW0pwT9LNL2//WEtuC6lef8Z5WasUrQiCWY2A3rR342xcCi7s9JMcgQwXHHtySI1Wk6vF+t0UG
NYppwAOvjsAiskc0QW1Np3WVQs6C+83eooRj8r5u9gGO6Db5zTAKmnVxAUHtb3GqG1p2TcZQVO9B
ReXdMOw5NilEMBuEF5s=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KVls+Vi1daoo6gixacoGC+YlExJBhqU6fWZiLu2vR7AOcRFGZrc9vz4Wrb13xk91ZxPYgqKhuVEC
YGIeRxZsehR3ZVlY0OelFP0EcFpPI3yklZ4pmPyWMMrZian4rdVsRQxiUIfr52oJ/mlN60hX8lqh
vMKIVv8s8LjadpJapOaJ27OclTha4o5Wg7+JatGvZ6S6o2yqpITNhs3EG6nFDCvP9o6YS0btXrMa
6RIIyzsIJrzf1wek0CqT3+8xdYczxEjx+tuxp5YcBx78Hq6e0TPoqTIG+RnSorNphvjMv7P/RdvA
8qKJCysBBrJOjq/XqLGtIPvKIljZztx6qk7Eyw==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 32336)
`pragma protect data_block
95MXtDrRh5KBGuzbCwB6b1/Td3yWNApr8ktGA4U+v+5ykL6UihfLHCs5s/CCRjo4baT9Fp3S8le0
U3DhaiCEeKspnqbi5+G0jV9mvvvMYeQtTDNebz/3EI3jZA2o31pvv1IzBgBvS6M6cahzO4dX88jQ
7q7YO1+8T52doplry/2dq7o+rcodNt3gpMIlOrQF9LiyfJqy5yGpMGhmEGybCna/CLVgXmKk/i4o
N+z7PoByGVA11+/grf3rUjPTR7zNjLRUfEAMw6c5JucrSz+t7HvWi89DfS5Oss1N6+7c3DNU/Wyj
XAw8QE3/5UFuT2JkcWXXELlr3CC4SFNRIAx9qi4exO0goXNudRXEuMjgaRcuwk4DFDY/kiNPOc6Q
C/m/esb+QnRVBza0SuLKNAuPSzZZDC/AC2B7okgoz5fddobZk5G1d1lnLuf8mJlnTBT5OxrmKqWT
ckEDoH9L9x0Qi5xzLoFPYKj49wbskn/eZNve9MWO2OSOBD1eDj1WTAa03JmQUWwRVl/DXwMzLMRZ
SfXpsi9Rk/94pfiZ4O+YtqkZKJY7OCegcpraaYsvTjx5rJkLedb0sSUSl7d83Irzg3gxjgtGCIqN
iTGM/BLyMCN3ELvojl7EhGpcKTJEMJZPB9WamuhtxcvHbR7O5IVjhd+ymFRqp2YSZvvTJtkWt6d0
BWzEedsl2bvvBWZ7D67hZg2/sk+oP758FI0HT25rfIgcAMvDneu97VZAC0UwEpt3eo6u4DIqqlah
WHd9WWJI2GGnkznx9PowJ20QsMiU135tjpqmotiOCUTwIUCxhw5RVHUkyFn+ufL2siKdcnmmNeUQ
9peSRB8V5/zwRy6pI+SrCIqx0aPxy05Tz25yxVWS+KPtg9inFvlIDxdISspzAntcU9ECrcKroqsu
zKNqZMRfOD9DjiGBthfgSC/6nvokS8RWk5ivIr0Oaio8HaSrSmOALMyXlMi6x0bZmpO9iKvgOYJ7
1Vko/rHmRL2tVassustpJ/s2Z41uponRLwvTNWgGeCr+2V7gWqZHZdhdgklp9jqWYklgu1oTvS38
Bn12oVbsZEEM+FfDlEwmBnpvtKsB40nRwRu8hQlLp1r9/qTv10smByiZPJKCEiwu/sms9BPgNaof
eZMSSKwZXTKq1n3Wddaour9CzP4EE7Jf47VwXDnGtdT53vxD/sIRQ4dPAGc3V40WlCgfUEiBF1yd
aDdSXFN63jdLHCZQtHw/4z06zyRb3Okto4ACOJ8uoIiipx01+mBXYQP/QocxtqFPXmRdPg/x3Gir
act+ok5lByf1eKx4d1rHw0TnEOkUt6/s0G6Am3LY4uxZ8YrsPns6ENonXQpCbwQo6vBPe0ROdmna
4Z8CYgOkx2+6aT8UL/0YkUM7Him+mNMKTH1E7vovEIYouNDOz0i18fRxQyxPOSxsdBGKbA15BLJ3
KzHJaXmjuCeKisxonLLAyvq2aU6DsFhM35jP7OfbEy+Uv12YUWjNcAgKfP7W5p0orGCtZ77zs8RR
z9vUbCItx0OjLCJERgvHuvhWnNN1LTn9wdPvDRS+ZcjDNxgK3sQkPrPWWRtuO/7RDe4dBRS/GWpm
NXiE3KgydBA1EK9cvvuBPhWuBSrvVgUUpL0Fn6H5Q6DQKfWTmscePtHEp20z0iGJcHccwIk+GvDX
cZYRby8jYqJDklRhPJMfR2HugTvb4nKBtJ2twPinCZUVClfS+qYE+7dE0LftF7GW4ab3EKQ8zwie
pYRfHA4l8FkFT8WjPJKYpoRY5r9uDs1L4UP0+NslTWHnMqQV2Lyr1oUqU/ktZPe0brihtfazdQPC
5w8cpcQOhq0jrI5gGtZY2RjKqVuMFWSz4FuuTmjXP3Upxl2H+NS1bsUoghhvnVfselbvrya5lqza
TBw7h31BIzj9Oko7dkprtZpGwgTzkm0XcxgNsygrjzh3WWoXHfO30v+XEzGWyc0M1tK7Tfv8UiCN
P06NjJhUbVhRR09J5wVmEEPoZtxLSFnbMz/pOZkl3tl02H75QNfHw4/OBePIKm+z593UhiJQhW8c
C9N8CgTbyNyV/J376h+g/Oh2GVK4hic3ECe372aFp0ThZLERkd43JzZ3pQckPJWvWJuv2MdYbtho
Pp85AsXoE3KlBvjjoFOnDqDRH++/5eF6MUEwL8H4agNrtU6+9QHzCFVGhqgeckxo7ErRmXO+aWzr
dtFjtd804Q1bFvk2lNnOo5Xz3KGQRd27JjQL7LpQrJghriaEblx75ipJAHOWF2BgiBK+nW2KFQ/5
xF2wKQ+N5JagdMGWiincAr7i1DVF1PEM7amea3AUTGhWbO7OgZq19+ggvzPp8HZWXL5NCRF9dZsn
dk4ZnfjVUV1IV/n87A4F72oubopdLFKTD/d+Iqa/MYHAj+V3WzadGFQLir2AufUDRo8vH7lK7u7i
SH3ujpREb8LmQ9DjlRJv8RV+VZw+s5D/GFYuTV5Bnxh7MLbg7tBKHB5ltFiDZcXMC6nUQIqt1bL5
38UeUAu70SagZ2ggpErNWaG0qcK4zRzwkc1I96ZgXcQ72xAA6xvUFgZ0VDGM9ZSkXtqoprXzs2oR
ietA6BaBKmD0iZtEQyJLF95GIfqEd9Y02CfohUl00hHwwtGXmw2Q1tNMSxafDqIEFuxEgP7YVR8P
X4FQwjSNnziLaVJ1TvitJ7ReJl+5IpAJsjVYVpQFLHqYqsy1Fz18M/fltzc5Xppo9VtHFxE0W7MU
3DbVKr+HZRJxy0+vVlJU59868YN1IGPwD7ARV+cOrUiyoT3msoL8/8m4/7+eb8v/B9mzTM6JKi0b
zXSPTYMKsYeFTb13elI8nqHf39HRDPa9tf7RBW2y/K+VPPEd2PlXJ/6iaWXudVtRfa98baWCUSoC
I13zmPeINqqteJ2GDe5nlcJ8UIVj+QnxPW6BCVd/BtT72E0gferFajr8DQsu0ggYQpMCDbb2FZu1
n1YLVSNHNEZOg1NGzcxYjQ8J2/ha/OdYEuVETKd751nRSSg4t/JsI7v4/5fV66tZfviURG6iZV1L
tPfm6Q4BG/Zzb/1sOzpfdq6PO60vFcBY1P2YG/rvR2Y5z45BlLo3DkBt8WIHwnKE7+7FTeCBdRZS
yWCCTe0tglH6qniezDJ0AA89qizaQYsI+q3C4EGnm1qdkTJbGkFwi+9Y1QDODjQrTYFNOie8fLyD
4A+vVhxJG2tCmCW2HcWFK8MY3U8sru7LoDXC71sLdEhDT7Fm2aj/KS1vCLgTGYrcOzfBh8VoOu6X
9ZmWl8p9ql1yT+qutjGxy6GfrjxKK8kA8MQKgGoXb29dKql0vPxWj/9yKrwKYi3UD8Wlg8mSzuFX
pIVbtCMLFSa2+KAm14RlewoHz5810ut7CWzG7tAOSH0shDzaC5FuowG8oBJ8ItBUbjEl1ubAM0Vj
JDaO2K78M4aMVfg99Ya94vzSYmIJiGNh4iUjRjUk39Ie50sU1t99V7Zk2yjGXHr+oqVVXJqD2isH
nC2j7cmfJ3QD5hfqv57qjSJJEMbWRpTvKc1agaR2YiO2TPb+0EBWV+/S2aRdvViHWV5xLBhnfSqQ
ZjPEWIHHSWe3expg1LGQHcetAU/BsBAY6/xdmQIn+Lvirq/m8vKIaP1OZy09jHHD+y8QPq1sjgfZ
AewpHxVoImsIlE8nVXe+F7KMjmif+oXDlGOBytKuFyVj9SHEvpEYW3bfF4e/b8nxZPzcu5SxL/XM
PbfQ0ejS4JN7FebD6LdiEDH2Qro8Xs5QH6rkdDtgD5yxYFvXES7vqvYOIaUZZrrNYDVLqprLxyUf
epVD4P5zpvKXCPy1jaEjM/KnR3MnZxWfY3ERQhVj8RbO0WSoEtKhg2xfDQtBYd4AkiWwXTEEPwtF
E86U8m5jmOuBHbjhfsDmujdvrjPTQ890WUKkmOV22FVndAjyhtnohcIqOWyDcPIztUOHhpFGkGD4
GN8BNdbxOjmW3Ou5pg08G6oxrYl1wPirvJzFfBtB+L/unuUzej85COMitjjxNti/j7lLEV2ahKXP
LPb02DSalVCmr4d4S6Y6Jk7+X2KsKke/kyXyr6E4fU1ceAX3s0s5BgtZJh+lY+6gqim17UfXRTWA
/oZ1437H6S2+d0biUO1w/mLGa2BZRHQYlx8ZfytHMgLKW/8MB4cK68F4c0gF9ul2jiqyCAo68Fh/
mLlHzagzB0Gtt7TCl3QoFqLYil9G3HUWxONB8KRAdJpe0s6liBNpbqJwInGdmZFWh9tr8baWZTej
2EGzbI6Fu0yPBH/DgQaa1T0nuRN2PIIbBgeri043xqlOyXGwb4bzIlm9KVQtYDdkfICUbKhWZYWV
+99XUQI4BDRG5SpJkaqyqRL09vuSrIRZ2yhNAd/5tE4ZPaCDfknIYF8sIrjsyd+MsfHqgG6IbExj
p5d2fZFuI7a8UaTwawIUrpeFkK6VqtLvT44E9ovgPmnuhLFs/K0nKB8upi6EuoycSbVAH7r8pNwy
DfOAMy92TmHfYW4JjxfOxIfGARgNvWTcGXyKSEcNWLZRWtdBmNkw1lLsJPhxJi53Rtz8+xF5CiUP
NCzKZacU0GxfJ+ndkV5H9MgiARzOqzeQckvBZPp2fgzrPeVHsZRTxnTdWFheMD9zkGUljUTdBpWd
700yyoJkh7d6s43IT8ufth8KBBtH8uZZg8Jsckqr276JXSakovl9ojbmLYfuo9iJJwObnhoaXA2h
Xz+f9cymLM3GjFIy0aYQdBWNyzfD7db64B1vuo6Ln8sKjzb0ncBo6gE2njtmg8dfMvEYbzBB5tGG
52+hh3JIrb8DL10Vb56+pLiahQch1014JA/MFthHZqGeHwxTUet6C+dQlxXB4QQ3Pv1aF5hob6Zq
y88coATIUPoO2YRfZwl3RK+vPAk5xJ1h6w/MFIWgfsxO/OzNzdGXlYozVLIDzvrsTIYKwpyeLADT
WNpnA8loi8Ji6JUUnnIg1oBJX2efhxvHWaADkmEmkfkaDoYF7vWdkYFK0Ddz/DgL/1/r/34o1DUT
FsjJGmtxaX8UFj8eJ5T652cisM7EcK6NPTwfFsoMZIIVT7vu4X/XaaikJsPf7M9FCUcQ6BliRRlt
t+sBoABqfzjksfTrRPzgNZ8Xnt6QGvz7W1OEd0LdD1ukh0smMdV8S+607gX10yCch6l0winieJr9
FI6bxENdl3AR+/jafT5zJzO98hiZxW4eUqfIpyfrT2XbftumsPoUt64oYw7IFoT9HnVSFru5E9kj
8y/chEFRRzq1VdL4IZZYsO/kT9z/osxHvTygGQZGgUx86z/cKVYg2Axg+Kgdw+L5iwMx/ffgHXR1
MZ52XGkrFDnuW5BQtR13Tw3HPg+Bs95TtUlXkRd6nQRPtq0t1px48vY4eiKUozOcK/Njufvc0HD+
iCW4e7lq/flOdpNUNnjZKoYRzQKGPsQODI2InixW4zONxOopg4YS59uMslwGbODhmb2nbf2b0pLY
nxlX4NU1Hmjw7kh6PUGRIjT3+qKK9XKsKWh7BHZqZwlKTxEiDusA77vOTzokPNJOqu/+25MBDQI1
uvHK5oScebAUym7JK+BSMhL2j9Fu2GZFe95aKBPlm4yP1qc7O8lRpWX9xI0Clco7ffGfsT/zUeCp
dgpZabhMLSA0NL71MbmZCAvxCJt/ZFNwzB0xiIYlb39uqMqMPOYoom1NfhsuFP5qWXVVQRctDVzx
g2ay01+w3LZLrXV9o83rcFCrOQyK7TV5gu+fC6ajUoY6obalG122Hpk4O9O5Hz8syXeEhSYPwCPn
ZW6TnBHcw5HUymVPdEg1H95jn/QelT75b9P691LO/+jY3ZhKC9sj3Qvh0yL2ECLQ11WPDwDgn46o
Yxu3w5oXm9CTR+m8VCGLCMCaxmRjBt1eO9/Ws1zLaKmEoHUIZRFtPEqSZ9X07mRLmC/BkcFp7HSh
bWQfDxFU8Kl4tw7KcS8mrBenFKPIMEXVNi5QCE5g7Um0vzFcnWYetMDYeXRTR6yBgxn/pIutZz7H
ZT8rG5zrDPmgfr0GGh9xlpT4558qvJqU+Y0LY37L7byN+/Iij4FoOSlFL2ukOE/a9XtZdVpl85x0
UiX9LtgzNdyttdDNdqj/aOvLygOnBk6vDs/kKycmQPfvgHkH7YMWIFBmNb6EvhnDFz5MIERemfmn
GT6peSTqF7L9jNv4BKoN3ZwGgKRzuV5iuUtBK/71bg1vN5pudeRjC+l+Lr2VDKglOTx+LVgtFDS/
UWY2LXb2D08uVTqie1hr4IiSXYtFJqHYxok1zC5Bu+ehGcnlhZgLohwv67BTy8y1nm3qOmOwE5Dk
OU0nU4IGWcCK3w729iae3a+fKrw0v02EslUFbi9xbvvBxLtpa6fs6tP+WAxAR1FUe8x/RDUAa3C4
rs2bWhVL7PN8g40t3tryUk0jt/MYVT1kneOt6yS36DWUsqUPrSvPzuq7jSdtafu3OvEeBCBpdDKy
DXk/VTrkHfc83jGHt+CgLSqBoGKAzrqsKQeVOMVTWYgLs70a4rzaLJoH+x5668oHa27l/npC3TIX
tu4vLF9AWLYeFhH0Vk+dzdKP43yMjwLYAg/Q1om+1IrZVJ0ZGV/ZApEP3UBQeF0aIqeO2hC1vj66
kVqpYdjZleImQEaB3hPAZdCs8j3qnrS6MkrJlSQpgmyQY4bXLRpLUwoGefWGn4H4llsPCQQdcMnk
6bhHa1uE9sZNbyvauXSyFl3l4+foOrZ65UrqVJk7ce6SAYMrrzxpwVBNj5K5AGzk8d53Y9UWsJ3a
IgCM7K0mbJBtCK2iyF+8U7t1xR1ZthZhR/HIxDtv/KWJ/1cpvA8+dLJJyXqSgaXK9dphfmtMASoP
qOfuSEiJ3LNvWXCIMKH9xE14FMTimLgOvhVkGsehezZkoVJqWYxPv0FcylgD0A4wV6IELk48dFYU
cgNCo28EjDZklEBYY+hY/yx/dvDqsTN7eqPi1jN5NpvYo57rhjidWz7LGOeuuJvOXD7TRKEJ4IPp
vHftpEtMvaQ2QAhwmzAk8xJvMkog+IuDPgqYRZUfaYCbgsP8znrgFqN3+7aAMpzmMy2RwOnTaHAt
UDfLlfnki6elgya+xamsDde7zEU53y330XRoa1GuLAMs9aFWSiEYaTinNmSxNzKqXHItRB4fsNYR
TnauMgdMXMO8qITI9VKPZn19SmDBH4fzpNFd3Kw23/7zC+hQY3z9HmUyKGkL2KexGPlNTWzeZ41x
YgNTRHu3b2QfosZVKkBY8GEGSdr4Obf0mnxnBVBIecuYFb0ykF86WvZ7Ve/6Ridq561uO8Dl2/K/
IFN2f9oFDD17uf+CmGfFojLoghF16RtD+mopgUsfxCnet19Pd7cgMuKYwnaFr+MCp7v6/RqfsPFU
5s8JuFeRfNjgOLHmvaW2RsCXBD6WrruAKDCJr87spb05TR8ygLtzTGMsKizK9Ub22y1K/TvzmgXz
UDthtLRV8+obAm6EQncs9t2N/lksSnjxGZsm1VNwceCI0vXr/012xQvtBp0mLO5J18N0/g8oS7uV
+PzWiwfmlu8BN26Jy3H8DN8PX9uKmTMgh8dDypjpBVZAexnyp0vi7amjmGhIdBYzzRyVnX5JESey
d4qOcVyfK8Idtng2BLx7E+y3B4uOS/Yf/4dt13f4hxgaqYL8cSFUKPG8m432jJg5B0MqmsUw45nI
ZunrSqitBGAHTXq+Tsytzjts51nsu09/Z1YnAEUSqCh/qL+WclSpqJf52WkTVve7Wf59U7mUVy1x
b8FPNbHywONqxZETwPv7xRkLm5RLIP3b83STpBvkaZ/6ESbXxV1PHvJUR6KDsezzhroGuKVmJKRy
TI5TsEvYNFKd27QTY62ieb5x3UDyC2TUlK3AR4K+K1ODURPUJ1sHgbwJzDrdUFMfahffCM5Y5lQM
6y4dkrzgXKyF76roSZyH6cy+k6AnTyDM8/NLsDwmtf1GXtrfrjMaI4/OQHgrIlSu2Tkv4YDqahsm
k/7+FsuuhiFbHRYHDwm97JDToq4D7MD3YYlTHHfwvyZdS5tk3L2VNSOTHfHF117Ecww8SzXlWnH1
fFAwpI4lXwVisg31V6FVCgpfLrZLs+X6+m6+A1Ln6FOLJXyWc78kecaj4kXH17u+4+Yx8lpzMfLC
Vmi+GqBqvd3AbUuW6Yk0UyZgBHiT+nTT2rl7Md2R2spbYLWQuhzvoYDq4jmF1Hli4l5diLQ9+h8o
Odw9TebB48ZOxzM7PKYNxJlo462YdWLfFCbJMic/gScmMbySKCUGzCNtIHyH9l+b+g4hPTexDvWZ
LuiSWno1DdD+fGsi5gPa+FA+M8ZcndeTn4tqeaavD0yu4yeZkmDMzf4ts6bOrG28oDWSp7Dq23qQ
KTPfgtqKV5USo0DqK6JVMpQTIxeFYRJ8wwhqQiyqLW9vaPPQUp3I/WNj7uzhlPzvxwaEIaIG7VEl
GsB+jk/VQ6P/DgmZEE42Fh2BroTj3qyqmuJij8sseHJ7YYxiKzj8GGo7qSBpNBj71K8tFgUyAdB4
0/r0BnafE+xC/n4No25JT/pywUln1B5vyhSzXuVq68iRZuWk6oKAfntDha1XClMCzo+PXLstc/Dq
zmMr4h8r9OUmhDdyUhJ/TG6BrvsWslqTPS3YFD4QvJ9zSuGMHHI4fvFrScJUJu9Sce2m4PVK1Lv3
UbUPo4wOgdsIW0tvVAcjHJKGQwSDOruWPHQ543Gjol9D6eJplLWFco3n302v9Ib+0e2NQHa9MrlF
eYUarIyZWBvkQiZ2L3I7RkiW2DWtTXxYNBgE/nxga5XhS2SE9i3to0s8ZPLw4V6w7aAxjLaDwebz
A4N4iyIPd7KZWUxoBN20Jlj1w6mSXgg1imL3Nubx/i9X01jGpa7ddwqfra+Knmrwca1/rkHmPvM7
dq2e3tmeVm7jxmgJPbPtadSTkDymaoGTnVxLHHywS1DekFI/pw91FWCjYvwohfoXiMm4kvZUjOko
KVyhuU1oltS7PsX3mzNmwbub1G6hHu5pegK57e9O36jhyLm30Oc3HdGmz4gt/agcsEqYPAf9Sj5u
5G2DH3zdaUHQlaGzevagjv7NArlcTO7vQudEK6EwN1nMJw97sVpRT5YIv021FpGsG1T/2NBCZg/7
JCnR0DOKazDK0vV4O2wVrvFYbaFLTjzEfRZ8gCFG6EBl1UQusgPloJHo639Ix8by76sibkayT8X3
X2I8aqiKKh/G6rCakhGh9DaPXJuosPpdEujysajyv5LgGGRwiGSSV1UdFTxC/86/HUu5Zxp87bTc
9ello99p1xqG4a9wJxzc20+3xlF5Xr56599ceQChhBcSlLkT3ra3gn60QQEOjORTdysfNy27Wz1H
zjtjNugbY4CahPlprlrM+0O/aeOw5yzdPMuydRB+QelTyOK9eM6MHq/7ulVeoa2p53u/+gc3q0hj
FLdQ5DGxodgCm0ArMjDeY2qZ5YX5GfhWIui9UBdcomYCMe7R26ZoGtL/b9AuiKb8AJm2jEjsILN5
sVdPOOTbXIhRd5Zc1ZXBeLOOQXDA7Q2foFmpLm3sRWH58ZV8y0xd2k+KKpG2JUNm5wWfannOGFlM
2/bob8e9s9C7cC9aYApLzl3kh+neECrxLoyBLCyWncE/y2LCOoI008emi80jL+iVRrEx0Jy0x22b
q6THdSPctxD/CRGIfg7SYb4Gp7VPhK0WKjkmRlhmEZwLFhGM9ILoLJWjX0/NofJO5GD1nt3ovbb/
MmCMGbHZa4kzopFVBQvll5kKpycTmJQ3YTaQq0+/tul4dCQxzvq2E2mi3KY3jnf5/30czDVuEFPF
JwC4iAYEjqJQqULVyd1MUvRchJon87SUm2Ygp2DGGVy++Jy3u2gWWGM3gFtA9fGwgQIWlLc7RsAI
m98PRGecJSl1nR+YHuKywlbFnCESe3R3JtpdrILWBSL+vCvc+QorhqwoNNClEL3gOMEFpg6b+iY4
MmP485Q4C71pEIokeI0MyupfW47X+giEdgJvY9LDITJR0h+eJTTf/szjp4gTW4N11/aBpmpO88TA
wR5/8yRvzK3PEggazqGxhTYjWw3OJkQyoRBCS62uTGM1Qx6b4FnhPbJAse2mUxoFp7cY9lyq1daO
XXsYt7aF5OUhUNlSzuO1C0HMnWuZVwsQ8pEkpLmGfBXjoMqrryH5T5+wmGsZ1L5F5HPUB6igGqKX
WMpeLo/yX3GhaiCQNy8TdyQOOZorl0UyPOPhz6TSDav/FyE6ODKShScUArbOAK6gArLkewvFFQBd
NG+cnsFVCrDjb9TL0V3I04xIBRtlE8aXrSl3qiWQG/9ZFSyC9r5hAQjS4PZFGZpzVFGxBvauhqsb
yawP+fngBZ8nHnc7KOx7wqgIN2W2e6SJRDRYkAnaJfcGglpNQ4M6dPE7QMWoz7PZW7/j/PLsQDtI
lwtF3CtBEn4ne/cmgS2BMPtDeXImpT9ejBWadpctyNGuLWz2abyP3SJ2ZP6XjFX8OaAMaq2Y6Z6D
u70pHI0yp3yuGa7NvCeLYvNCIqe044J4PP/NinxeokC6EO2C4YkNncYpFL95twkYFXNPHMJzMvqB
o2F4AmMtgaVAF4sRgxjv01bJwmnZdvfmAHGY/0u5Bmfk79fnjXV4r4iu8tNJodhSTl2LWvgnlKkb
ZPyVDl7/+8p/M3x3pEdN0iNoRlI5pqym9Uh/ErKb+BAGcvvVcIELQ8HcYfPDBJQF106sK6K5fUgU
3/UnW2YrJG2MNc+yZCqy225Zv/RgEqNAMUzN61KPnW09IEgyfoXnYPPKHDs19Ica4p2kJ4rVoUMO
6ns/qxoiAp7+UqASWDd8a3lAA7CMkp8UbkZCJ0YEWhypko3HtWFeNGY4JkEGSt7SgR5E+g3aZ4NM
C/YZ+l0wUgkI+2CnZAaXGXm8ZMeXQVo1Ju/qszl3ju6DTsug7ytpXDhHlR8mxLV7mMc2dfJ7gau0
llQV7U1D6/BE8KfdDUsC8iWk0eAMM3owfT83CEnQYHQhh2GnR194k60PXFOkGsLjJU0mRmWNTTbD
ITL5dTA7TFHVS5HkRQPagP+bB0ol/8Yf1L3yM9T5nTvNH01sd5aTr0uC397KnLj25wRBik9um9pE
/+tjrHY6Gm3eeoOBtFt89TKJadAk5Bhj1ZNJHRK3Ak3FJ6o/GCfyYo1pyo0qjaALcLKmBr4zOQvM
mYod+pEYLIHUJz5XRvWlOeWyZrYO7CmMo/7EaeG8OzVtl03cEDK4yLwOP3x1r+8koNVB/u47E+xH
plXTuu9Rvg1GhMqTcSraayGYem8XzFS72Dn8FIrBVM9bkZ752tEFRwnKQteiCos9oYq22MavO4Ek
gQ5N1MwqcoxeUKxjClXLsBgzuZ406JMNFoW/EsvBHU7mbH4mXgv7DIXuZh40rO+omHeIvFSmPKG5
9L+N4Mu0UgWORJACNO8bDejPA3DNiUDq7S4+BQfsal+Y+vIBVV3tw4yDFiCwufXeMxvR7+Qr+1vj
lY/9seJY2j3wl/dIUpEjVt7iuN3t7gYF3MMMtkWMun1zSp2z53e0MkNLoqqBkEYiP8ZoF1KvDBwU
9dlaceVwVdqC2bGEfqQ9IAJ7QLy8aj5GY0YSK6Mb6lofHUtmiijDMKTTaKusdl9QCa8/9Ca+81A0
mHJeJnVgM5U+cN6XQ5ObhIF8Xoj3ZR5ALxh9/OP1c5e9RB0yVlqoxRZSZR5cJBClwh49GCOASRoi
6uVxwdkYQKB4GV+vHIdZcmV6E6bY9CIonc2826Ucl5XtisPVhchYNghjGjn93HFVfxsfytn1VG3n
NNrZs/xVGwZ2DR5Vr8A2KjZxluCPGBK6zcwmVRO2TYAG4Mk6rU5E+DuzY928OySuKnnEpMJIhAqz
kaN9r7IRXGVRvH/BqOORrAcubd61ZWIr8OObEjFhT9gs3LoJ1po6CjVvsGGG7FhaeOLJHtzh3izx
Xv1o1VIuxCq/bdg7qnjDh6CiATEm3+nfbsCtIyV3mDeUZq15dvNiCjmwdC4hfgYiAP+LPQZ88YOp
iG2M2zv9+14wOVrcDzikB7GheodkH6l0nKIyFm+PwdGh99CvuGrRW+8AW0h4TMZ0cxd4AReXkB+B
W9Kn0VIEos0UKGu8U0nug/qmbn2iuOLLTOlmAkyabNbeyNQpUHkv91KdaHxvcDA0/gCFLTFBi4jm
eDip7YpsX5x2P7eQKF7V0KHenhz6nCvCgrwkP5nruEthrSTv1L70q++GA1fIjkToH1CUTFtJROE5
rLwZxkGgqgSqctl9gA8IVRE+kRLDfo+gOLCtE7qTZtM3d/9dI4f7J3YHZsKE/bc38WPtPyFOETqk
UE2iar/S2GFPkfDG2QNb/LSRWej5pde3+PFZce2kGGjXlv/OEAxXt3bu9EvpvEYUnEVjo0gst9nx
XbYVP8SS28nKA1egmysBnr72fNT2KdVsNfyjjU8GsNQRGlVlCzo9OAy8Qdup8bFEhJaprkZ/gnJF
p/EeLCI2Yb1Gcy4zsQM3v3g7uvkrZsIvOE/lb8Yf/qW/NUPGcu0WZD3GQay8O8MiKGbtTHatY7Ud
Vjt4oIqzusCKBoTBR7xnp2T3zoG+FRJ+TJVsYVVeZECNMeuR5aoGJy3GEdnC/aPVPKYX+evf6S6c
upT0q78X58X3JJFR/VkZEbwrnimsjGQrUrNEYU4xuYUEeIiNOy6pSjw8BquH3BAuNdoZgqZWDkIP
4kcd6jmL6TjZOPiGde3+0YfxT6BG0nsWjy+rjpCJjJr/TVm4kdGLvXyqIaqNjKNY8yCHf1KycLnQ
7KNkDrIPWAz5RgYn/wPqxfway6SQxf9PaU2BRpYxI6lA6mqIwFVF3jq5RZ7NFVd2wIPOvvd41sep
i+x8AnxCdd9PTXbopKxSAYqpfl9vTpuplcRL9CPrXVFDK5LSzp7euCnyA3/0eXWReJ1uKL91jNYu
EamiOkHeFJvB3niQSvFgT5EJ1u6TP/LfEwRqQM2ABlPLIuiVYjEIPAe2DuWUKSKAbJsP96QqlLES
1fhGI98lG0iv8uNR8lHw9nJmC7FGNFuwelvWbPXfw8bfFbXkFeDwtK3w3zgfXRM5AaK8Vg3jvu1y
N8DKXTWilSsLTgLr3C8GvvtAMunRweer7yp0H7l5L9cqTU9OrFfxLrV7YS1JRTwNfR61YgpoH2/W
3SoSmzoyzxEdM7sK7FU9k90Tifg6AnStTT0HYkoTRLLcIu/QYkD7vg1D9ookeU2iYtsHVmyTopbQ
A16kI6iTa9X/RIbgIEcVH5iF5+nWgGSW28l2bsyqPYbonFQhM2n5u12Y97G9MaVxTelyiLQ9pWjk
31WqYOxUbM9k4lYTWwLuPNjPybZY2xu0MSa6LyodVVG/Btgo7RaGeX3KIRkRxNbEDYIJiDwqGffC
7KPlKOc2zHevb5BnT7t6yCJwtWG7bJ0Fe5cD3qy3jBmgJ6oi8XNbeW6Om7974VfeEY2H+RYNXKvg
PU1qSk50M1gqkNSOmOBElyIEgVdR86cbLvPmzRmojMgFhelL7CIaIdN3/bU5LPb3hlKJ3634K3wn
8Yd73LQh8akFvTWyeb0Uzq6E/6yWZdruud2kWP6I8gJEsx3i1elDNcQd//PkBaLCaEPtvMJfxroK
gf0sRg5i6Pqd2BZt1oi+nzbftO4hkoJrgFfPWdI/4dejrHlDMVamugpHlKWk1c08XMOcG0byeGl7
RyGGHML6u4vUHcmu9OIaVPTLwrCeboEFCwdOPKuuM5FwXWQWjww12re8nvtaOcvMDV0LFtEX7jET
r9I++1//N6dvcZDpLReunex+7oIIfN3o8FF+YPZOPCbWJyppvd7Gu+aSsSQEmtmz5hhAJqFlncSZ
u6a8qJAPYrXAEKfvYVmuEi8KY/z9/YEjGQN6b0vvFgce2giLG+HY0yp/s+dtL0ZE1VZl94AUfjCN
i/c90+3wTB15+Jyq6FtPb4MrpZ86kyzGRs4mniFTFl7YRyR/PaURrB+B07LoUWqBWSgZig6Cu0KO
bM0KzLo7qt8locK89mlL6L3tt+1LsftJ6yodufKOTDyuVMo71nVS5t/Ly36CLwGGx3TOyBAjU5mI
92VEgcqagg8QRFrUOtv/BAxojUgfyg6iRvLnqFXhdn7XTLgmhc8ARWv8tw4fQkdJ1Lu3H6J1+FVc
g65OEYb+O1gOeJ5+cdLRvRmzE+2ZwAd8iZZRhu7gRhP26058lqYLZCgWjcAkL16nAIiBb+7pVkl9
V7qQY7/HDe0BNIUd2Wtf/ZgnLoxGTiGzm0Jp+x6MBnLUr1DPq7jQij1T57Lh9mpOFFG4MQO0FSOm
8JjWgdcvPS4boDaOD9zfSAHsOht6yEHxf0UmHste+ZbX31SLY/+MwFQqfCSq6iGQuekhgsMjsXyV
fcVgU0ErtgRleCh4BsSbK+G//8jHzCgFnvb2oK1yy6EWH+xQzTjzh0tOmLTbNlYCKGVpor4uFgGk
e2hbupOHi4Tcb3UI2odLMABLaEsNlnil2vFXRTvmQOpA8z5hPDKp9tGrfjaEOEbUi1c/S3maHDXv
F9zTN2AV3i6O1p8o5OzO1CXl63fokAaHKHiYZaiYe5fqdQKJ33I2Ptkdyyq15iNICecrom6I4SXN
18S39hVAqLw94ZWyOgtCnmUkkcJBxrhk1w1aCFO1B6/MoPYVhmsn9vpAnYa5FQJixgFJ05d5cfSI
Hc1+MPh4OytscLTofP9plFIkpk6W/QjzA8Yob2tV8cUsiST/ASGGRkpLc3e1uDBo9o6rfyeoXsyH
YM4JSL2jzm0h5OLZdipq3Jbkfy/WiwPAmX3MOccO8Z6cXA36hkp6FrItsnqGSe2buWQ3LS7bHqB0
5aCdzmGlX/4sQ6EBw7FcLNE2jgtzLNduNswboPrJ3vuDl6z+zVBuRxOVYPFrxCOsNGKd/rvuEXdh
GRDvyfPiCmDcR51zFuwlomMudRTERkrcipS+Sz3gWBsTzb0R6TFEkuwvtxXV8jPEKaq7d5J5RRu1
xjfp/k23KIcb+TYmYssNGL7Mzqe0MuftfEeTMYdjN66TIP3/Iw5//V1cniu8ZKz7rCe1wNtD63MQ
40DER2q+GgrSpFdmMdkpIXOGoYBcrTwk6W4sXi5EB46oLUe3zGvmIE3mn/2Z+iFMoQk148+FWo4b
7WW1KeldhPBCiSTY9eWumPONrD3sh+XgnUD0IYxpA8T3aKLkgx+nowXJVksNqBF6/7n/O1DPZhYk
Rjv7pG14gcJF/9X4c04hYFOuVTQiyM89T84H77mAaq4uDX6ewoHmPpw8xKpYORiAq+auHtVjgpqk
IZ3hhfYt+LVsD/dIqfrWAPZ77Dak0CHHD/qVzUbjJyvlqvIaqxbqN/lRDVzrCSFv1GIF/O/RMsP9
r3pyiFKTede9pchRn2l1OxXGIKSQVHkdg2KetbZJlGuE0zStq7mNLz3R6xo82+TL03FbE3q1LL57
F1VgOPLaPXktEOxGRKuRt0gvDt90H6pS/OCPSDW0gkSBcrYfFRWNwlvR42QpMpUNticy0QOKkEmB
DTI0+pTqvAjGjBw5gCzTRztIYioVbtoIDQ1PqIC1cUfT7AFnHbtNIQ/F5EG6y9a8TNSKAv2ZBZmN
Y3EXoe8yhSKxwkv/IMYQUVJ2LkB9V8Y5Qrj7qITBngpvwCmcbItwBLgbdJnHkKqxrfAXsqTsmyn2
Kpv6Wtb3iq4PI8FwNLIDPN87c38wBfx7wxPzQ/xt8JhwYAT08wwsnluqvbboegS2TDNR6Du1H8UQ
T5hCSOBC4LbUCn8jrI1ePQ20ygKJV+lmtPWHbGwbtKJFIo59Kx1kxUTMz5/M5y47tXVGNvW2BBxr
B23Z9OqE1L6hpyhCOV8kdaXhb+JgzqEEJZCqmjBbB24kt5Xuh9k+Jo05kdLSJ4WxeUtrewDG+QJB
Sc4kch40VxZBLiOrWMhbazz0ThD/dBI/uz8u/BM666H7FgmYbs4wkIKGmSydx1FbJl9JqMb30sRi
mM0vMTLboiTgyOdumQlqhrd0mRI+p5CdLnw1uo5zLkD9lrmVPwsciQxPzU1G/0UWLi6fqB7dM/OS
h42UwNUP6L7nF5hJjkrlY8BZQQ9q8wUekRbN38JrLOYVdq7U6BC+JCPnaPqK4gNzbvBiqZ9kkxwl
tKub+8aw9udms6tc75W9nUgt9N+8KddVfpkY+Mj7SiHzEVY9sAYGSD46C/tnRk9gF34f+A7PXTl6
aVBrvK0WlN33hQOTUpwFNc5VU/4+IBRsQx7Ki5WS3LwrHgl1ZuESoSM+gfMUSO2Sc3yfeZI9EWdO
vjA5gjvlin6hG/bT/V/+NtvFg1JL9JMGzw2V3blpFG34adKlgTX8e5JSEKE4k3ElBH+q3sAEe6aM
jQ2bJyE+WorwDh3TX9iinWsVdG9VLObYlB6hFY4+QJPUtfr9Sede4tkvAD0/VfRi6kU47XM6sDdD
FqTcZ+SsW5D+qAsfGcb8SRuLb+BFn/rRjqpLBj9ScKsbljsTw9uZr44HntBhwfGxPJQ73t++D5J8
ZDnk23JFKvIMlOogLyO+wpLyNkCNxzxeToAsxbLhJtQnIEWyctVXSIchGqQS1tOcHsRlF7NvFNdn
11cMMa3aO55AFhNL58lIqecoWv+FB5w+Y9/t4Ip2yiv+F1oJTNkRobi7+ptQFoH9czBhFn5nCWWP
9EwlLldr4OBnDY+iZW7RiTSnNGYAjHK7R3omlb+4nPvkQVtpuF6U+tFmFS3q2eWh1E9BfLfK3Le4
BUaEZRJCHiP5cT/VXnsUeUOn9Nysh6r0A9isxbQQQs0DpHgUaX7XVXqPu+C1XOjp8++L9A6J4pwg
W3cnw2z6AGOaRJdgZjqJjiytHmuP8O4+FB8ItpCIpFkW5D9V3e/ilfKyn0hXyQOSQPhtmTKbqFw1
iW6FMk8qdfyWV+/nl5g98ih9JpqIQTHHBrGzA7r/29dVS7up+VMHrog6FK7XnbJTr94K+uRYlc8J
TlezoYc2q6IfO7yPMixYBc1Wi75Dv2UELhzkEfNJsbaGjCTPHiAdSQE8yE81p0E9LNC35i/8pKep
vJnLALkY3xzLrADlwcYUvXicm+XUhpRjDiOjGzX1BRa2OYo3qGhS2GPKhwDH/rRC2+NvXikU9waf
3QT71bLRU/5MAsXu3/ABJlVu6kExwTsSSzWLwTs2Y71LSFuHnveLowPzzPnJRIhHC6qR3kSFgNGf
KZ7YKhYLCGyYL73uvS0AFG9HVz3zjctmDzwFgdb5JxJcdDvPw4RYpeIrE7dgvuuVoon2aDRO/y8D
fpKyGq2/EtUpZtugEx4JUetFI661Ppb2/HHhlrXru3ctlYuJ53i+qJzckKNk69hSqnzLmmpHW/MH
bQrCOkmA2Hr3Une7IrT4qVdHuvNqBrU/atcZHr/qzLR5ajWsow5+QN7eelnMogUnL2aPswoeDG+4
4wFVqxdNq+xxvu1a3aM4np40ViDraLEN7hv+4TgbMSH1gL3mM/DtyDSm3edncbLr7c42eFMABzsI
9gyooKVSLHvo22/34XIfwg6GpNIgquSXOUoMI4Wxtl4L9Jub2Uge8Vm+ucNXoU9/ottv62+e3dDJ
ZKmxkt4u3NoCdgUOV6p33JsbMrjgSdT6JtIRNiGIvJuwVlRb5hC8fklmx7pZFvl02J08RqYieWYW
c9msbIOCS8QFptv+hUcZl/M8UMCV9JDombvMV2TyVTtsBe3+HL88JxNNy197fwllpgmq7y1nPl31
CBtLQwgbE92wyHEoB2g/bJ3Ln8lZL/YVJST28oz9P59YEQOojCGkITKI14Yb/bGpD7uDHZfl+lI8
EXSZryWhnQs1LjLZwqxAo0q99QN+enUO3JULV++/s4c4VCpHF2TDl+J4RqVid8wcCZf7Em+ZvC+V
c6H94V7hCk6m9QW0jkU8kCxB3iHpjgwi/fg40mTOzzdEEwQzlMrSrFGk+HcTimo3/as9i5boQXJ9
wNwITLCDGu8Pxc6l0+13Jgq8PTozPsiqJFSA7zAQbQiX0eHW60nS1RR2QL2UB2OfprqJ0/RbFqcl
Eyfgufnd3sbyjZBep/HfyNAUaxq42FXl/EQToEUkfJEf7k5SgEEeYD0mkE962xGKFeUJ7jPawW/N
/GH2W+68xD6CbEwJ3X/KaBK7U/vdsDSu41HwHW9VgoQzqNb4rje1REmnM2Og4O28Skq9YSV4wWAH
l+MKuLqNnha6Cn7QNoAM/Y6kUIhib4DCv4zObT8bPPYeRyXxNodeHeUq5FKv+yIJcw1aSsWFsYK4
PDPC5niHy044zqICOx7PFyFpwrO9FGgTWjI1emDgNfJ4fsx12JdQYUkNixdBSsqkwMSO3Xnd9eqB
nR8q0/Q8J7XZJsOipAtrE4hVXDWWLi62TfKX50HtTSfUk/oc7vBX2qm3ZGEh5mVZJsPa2G7ilK9M
ninJum60BR1lw8AWHe2Fx7KQNhTgzI9D3qpT/pHN0UoIL8p8K67sg05eD6CSwt68emg+IQJMqeFh
+7BLmLaKtvPHBvSzlzwndRGcIz7NJfwU92Gnnuc/L1hp5KJq6wnnXA5HjyVxqe6LSJ9jOXfFmy1i
EzCDZYvKc4Bz7M/6tNNwfZ7Ll6YZsuUAy2/JKSog/GE4S/b/kXhZ7aaau8/0fFCW3GaxScflmDDd
zD401DbHmUiaLb0khEVG+B0X7L5rzLVq3AMeZdrt37kDJ9873jXCx2jsX2iNbAORO8OAYY15lqk9
dmilsFmE5NeQODryez/AW+lmyNZON1x9lyEpKsDjbq2EXOwOYEiS0lGKwUSDQqmy2lGaSi1Dd4x5
tIJ2Xc6ldlhAIDvE8wpC6j9YikvbSWOgbDQGDO8K79HwTMfTu1n5EgCEoV945iuJXEx7mlNnCnwq
rUUP/tI1LwS3dOng/rgRSxSwJCoCByw5f5pYxLHXbej4pO9fI2fCljuZ4wu9NP8b0+ZCw8f5ZBq9
dIDVHEIOx7ee8Xvu248092oilp6HvgtMCVrKnp1TRz9sGm7AteXXtvwSyE5euIrFC+CZTj5PqtvJ
IyLf9/PbepVGprT5ATt4+sARoAMZoTyxufN2e21xfOcgSqrRo4DKDFkOjnJgNMGoi0fbiU3r76Eu
rr+HlVB/kEEWDzM1BNL8NMoYmp6Ltnoeooe0d7nFn4eWXeYuk54gZpJJZC8deI2vu4QC4IpjSHR1
gUcxf1gqeT4TWyKSNdRHlQ6rjeaLaRByoXW6Z3V9gjYc1hpnpT9poX/ISziFbfYbDV0+4t080T7E
9a8lySKqEhi2Bs2JoYRJced91gVzGIU2//fjCbJ0OSCfGy2h+ziftuKv6LumsGWiyJMYtkuqVZsD
hP76gyTnNjU4cydmez+JcOW82E1QtMkJeNafswOWE8FlVRxyMjjzuT3gCa5vdCnJOIMHrk+Q1I3U
5yZxKqWRttrzIfn3nkYgPzXpIkI3cN71miDpseuxm7Gj3/FudAoNcALOfEIeePSaaGlQHAsi6dGD
zuUTZF60zEbgxmdErJ0LEBMKLAKir4TIMGWuLRkvWMdngBfGa74TF6jXLQCwnHAUXew7qH9S+E/0
xRbgFzVR+JokJD54TvjT2IM1pGUOO9fTDSX5d/lOgNi7owRqGZxVMnkvjYs3JAjxG2myigU2KN7Y
Mph0/wQ2+AFG4jLaaE1lC9wt5+zryzfWXg4EUQlTXTJnk0ODsIKm+L+L02zx98z9+qFjIPjonL4w
FaApgWbAsmSbxYxJ12H8n0L1gCVwev73AapspP9MxPRA4ztkFvHJkTzm6CYbJ07Myzwakz7XSGgP
AATxqK2apKsuaUehj4s4xORtpWqwKNZ+KkMgb1uZprA1Bmobu33DYrpEZ4s6fqsUQFVOk8Log7oG
s4QBijIum6OpQZK9p0WHCgxX30USN2hTAqE9G0Nip4kB+DSCDv2O7EekH8ud7MZs2Q323mPohR+b
/tg3CpF831yNWrBLzejNT4AG/mrFvGRFZAUTp5YGvk6e1rbmyJWsW6pD7A6YWQ/LI0kBtDbqf/zq
LOsa3IgTIfvGAoh/UbNvmLbvm/lNUQFAlvBnnJuvRZhMmkpC7dNmUFxnq2qnZCVlV3W/piUHmNo9
tr5lyKH5O5bQITd0+JzvYV4rvKKimDCAOEWj3s76YP9p+sln73+7lYmJBkBkJIA6VA5Yr/KJVeUz
y1msAByBbqjyHjNPA4ZE8EUQFQKcJAiPJMyPkDVRH/5Wlw6z7D03iniGjz5ZgXFj6Fds4OJXC1DM
awUPaAsmIK5NCCsp4AHAvd1dBUZBCbtvIsOgW/2j9dpIsr3jab8yqb/jfLZuF536UVNN8ivkHhhl
nkTnYKY6HucdlLvk9spLzubR0gD2hg3XBAT3CWyQcbikEK+93AJ8PFe9yW6WBHJwi/VvexsJUTfv
8/vFUW+3PRiEgkvZKDeQhlX9el4n7+dQ9VWyQULha4ktoFVwFZM1qPGJqphEXP1RcbxjLOqZtn3c
NllQ5nfGb4YVbWn8ONxSH9sUsG+rDKFv071oXWU+cRm1eZ6UbNKp1GQMmPynIx93s6D/nppWiouH
+DSxvl4PWpwoYj7yRsiFWIITYF4BwjfjS6xWflQVpddadrQ3prLDXBx3FfGHRNGDV+qh/BdpieM6
1s4xqMc129dHTY/7YzyE8iic+cS3ljpD/CbRBvFe1I6gODQKyyySpMddj2FtjYa/xOFtz6iwypjn
nAUrfqXYSfjsoUqFfirOMWRUPkXHgQTUU2tMd17W0V+lJRl5xrWm79xzCz/ARNKQ7y/cVdR4dfmK
7nPQD1wC19MX1DGcQMFa+ty1nMP6jzt1t1SWgazbCl6OIPTaHbeorPicxeGTuhsGaY0003Hbi2ms
iT24ciT8mAYz62m5OgkQjdF6/acjZ0ziMGzR2JDplMO1edy7RW6OjpjnC3qtIR8R8UbmXPlOz4dq
G1U4RlNp/H9HdXdOObqlco5lVAgMEonNQuhpcjfHqmBFTsLC9I2mRm1XezzBZj/hU/qDABdlsiQD
DLwOBS+pbrf7VKdGXFKrnZYGstGdADQnNvFAXIGl8m5whRSqJwVPE4qYn3kU96BGfM4A78mQuNF2
roD/f2H/7mixlXyadiCitEYgV9wd7387/sIzaU8DRzMMEVwg07tDg7fmpd61Rx7ceIzD6ECvHxkT
yhyNZ+BcF/R5Ba2csQg2Y9M2ne+u1M3hvIHli1JwGzImQjT9qvbZ36DAsJrUMMMnAOFrYysu96Qp
UuWdRkdAjYSLlVM+IYi4cTRR5m4cSNLJKHZpmEEq6wcXZwtaHICRnEDLd3XqwiQ2Qzd/42/l0TjR
kA/hXBQTPawwTOVOE7YRFm9yChZSht2vwybKwAZCqlNpgwKWp74UEoij2arT5nHnnlqkQ6ORwxr1
nUQTppSqCNG3N6capwqoJMvZGob9kSfWL8UBCSwa7y8ne1P9r33IaUP3R2vPtxzGoL1Cz5GXal3Y
qXPvXLcNAlhK9MFylRLJ5cxfjl3B5FV9EPCnI6inxhiFlDlzuAfdHoJNQ4rWnUcYY1Fz6ITtMkgK
weS9dMiz8DHTNTifnwxYiY7eOI2hvV13yaTHO4ZqpKJgIKObnIQEMoO6rppLxSpP1v1G61QW6yT2
XMDTudkX3Ct4y0O3tc0yH7zjj+ifkm4V+MeNwUnk+iIA0A98ZLl4yiD4xuADPCbV5WUu7mFlE0Qp
VQE97wPYYlb1zWGarVlWTp2bTxCv+EVAuK0oe+2pUEfQ36jtmKJ6hGfUo3F3Wn9ULNbSYar/ZOuK
7fPj3ZekhKbuF1JHbfs0VwOBF3wsNxe/1tprX7DwvYkwOJH1FVLwSDBcTPQRvn+/dBT4UiHzFe2B
AuBWeHvnjD1jK+BFlxjsUxTlt5C6bEzCt5vOmO9bGcNcOw0yvbi0sDTkj8OPvLlWzXUcQsCyxs5r
SoxRR8ASkEFpgzA765BkamgLoz4aFWG8wGuPewpczJ8XDLkC+jji9ZEKsQWn+kdsmItadEkhw/8F
g5uLiPC6Xkim/lf8CrlJWdbMY/7AGSNYiBW09/j0gnE2s4A15/RU65RtMXAzQNeG/5RN2FQcenvC
1bKtCpN1osI8d7NOXswpQUWHM/2fc8gInZo6pPHr1bD6bwmmBIFCFwKkZggtYwnVzDnAIK/sGA+q
H7EDNm+Ucs4+ny1a6TUBeTsqBvZx5/p7syByUjwx997Wc8IX/q9aEBJOhF7JMjP6fTw26+lXzxru
NfCz46oxGMcs/dabQ1dyi7MTTAKM+tYiFGZ6F2hoQWQpMm88/s1ehr2iRvBYHVSLvLRT59B7dRGy
cVEwDvkR4/x5StFhlv2CIKrLsdD91clf9sbOebPx5fQ7SZo1jKtbUyhUn5frDdVuLEvaGAZKRr0/
u+jj2u1FeSqJFZBe8ghiZ0SR9WN6vYioRQciv/pX9riXS7ruI/00wm0NfeNcDVCGmFmClzI3/i4d
d+AiXqhRVRlB2vxDt5lY5xlJXAojwtX19BtI6eVB4Eh9Fed0Ii45kQKmUSKeEAkga7VVqd4FLXWN
TgLcQIJXuokI8rmcAcvIrP1cJswgiotrreOdbkbaGr80yhH5ceBXtNDICegrDsqWHPVrde5oMWWC
PW/WZv1Wy43h7mliiZQB381FU3lHXuBP1oMWMPOSnz7+E3lANonRJYHufugyWPFpy7PTM8HcyCWs
hqh26vrEUjTcfyHguY374B3PBGttyrFOHQYWf6ZPqRY6nf/2oFLnW8p9pmmlOhJqhd+ow7jUy9gC
JEZY5oVFa013kbmuen3fYb255qQHlQO7O15WjWWqC0VIH/4rNda3R23ltDEw9u+k2+GZ1sYHJPHs
eOgRRCSwGhdT9DkVUOv51/OGrCe2pSwK1vIjTS9yhLsezijs/0gSUQ/nUytoBnF5tZdlSQzsocOm
hnExjTHg1knAkW9PfCmOKMok0eHA+vDh+OujNFtKF9bDh6u+wNBroay+a7xRjrQ8bfaF4ZKcwizw
mP65X/fl6tSIA4mYI/yFSeFloIzf6Q8QLQSb2UbHhueY+4/E48qS+N8J/7zGmnjTAOM2D12OyY5w
e6zdpeCTWh/+kPj8mdleHKEcns8aEo3vRjXTL/ryHUXQA/s14JcIfM935jIyOU5/PIS0vCdKOEib
Y4lul7qF93mqYDvBSDNAO6i9dCHNP5JI5yV4yg220yBoLcBUJCx5GugZjt2n9RtPA6aXWmULg9eH
TS4XME41kpuLEl7exVl/Hk+uSBPkNFXqRMT+1ifMwIdtuZLzbwC+3gk+VqqPpbDXdygRYdlrRmL4
T9e0ue8ml8WVQUGL4VRtJ2uE4XeOxM6PeE3CyaybR+WOhiwLjvmswiFT0T2fmX6PswniDxR7HeVd
vbkmpySFsn7aBTNiRHPMOn7fQtXc41giUiN7e5RkjPsDGMykv7999fHHng9n2eTwyV8mll+LPbvE
aQfF58a6Gv71UUjHet6egP3vEdcJ/o54HBDgz5VV91/ATmuMT30yX/fOOWxRiHdK56VMtE+qcMBj
AVcsjGmv3nK0JUxNzRPOKFNtb6UY16sslwZaFvItGrvldWw5bXtbZwbj/ZpRtwhldkWHBr57Gtl9
OkvU53TxQOL8bMStr05mPaDKg+Az21tKDQwercdx2H/O200CrKBlwqDWmPKTdWyyIADyyjUz31am
uLg9p1bbm07Prg8S8bOwP+dxOSh+37hi/5LeayVUQSCIhn8ZEvihei6CfURXrVje+m59kea0kAyX
WrM9KSe1C0u3DlHgDt3ED647iUWQgzUGh+m+et8xQ/VcysSEd1E68w9quxo34RRJtt7ENSXMAEVD
QD8bYFlhMUPQgLnfBL+j9CqBPy1qdAUVNJ9jB4Q2VxLrZGy5MkzmUVNKtT/iVw5qh6EaUPLiha4U
mnvyXFKKKCic4vwDQB0RyOEjucAysCe065Ag+oxMpey9Nvf7l/z5wePHpQKtgr9Lz0hIZaO0wqxM
tQTQW/lahutIBnp9WglWaphX4C3qNnGLGTKn7v6o7LU9UwDZxpNZnYxQxsqDbtw13ZF9T0I/yX4p
r2pptxY6RGTZYQNkSVzYMeeaFUmxkPlMvV1HOeyzKzyGfmMUYlvDXM7FOvoooHCbNYtgbChiStty
b43chX0XSjR3w8g6CWMpSzgCYXvq1MRbzah+ZBSCKfsLJtB62tp2XsHEfmh7u7uQrnlaEdm03R79
qIOgWxdjJX0uC5GGOPwBOWqUHr998jPhF7/Ya+MR+d8Tn7c2G01fsKoVxzoNgKeIol/Cp27+Jb9W
SXmjR1TtAnaNrpGDSwzvSlU3Wa+XlJi8tuBRRO0jATw1OxFg/n23vflAk76ez8iw29B3jGNkeigC
VgaNo7gz5Ki6C1JI99kJZxqt7pSHH9zLpmDBg7ofoL0ORewINRfOhfLTpFnBkfhhPRQRmuzKHzTZ
7+FRgpCAd0hk59pnCcxdnF2q3Uv+0CqTyuNnR57TsWjNXT09hkiafS1lH3KImxOaZFLjcLflAwOY
6oEvAvd33mqIL5grrS1oKBomBuG367Bx7t25Qrt6C27w5mfW7HUO5yIt8ndl9PduHHt7PWkCmuPk
uSSS8AlIkPlnby8FHWcBm04GBXyH/86nzWU1sd9FKeMX86Z8yi+w4yodXNFTYeVelJM5RaogRsPv
8tkcp0qUsw/tuRFoVNNlSBfHa43fVcJHp6f5247QoKQ8MDzyLvP2iWT+xa7MlK/EPqVjWDJr4VYA
vR4yKKl06pvcacN5mid9ouLHs7sRfgPBOddQr8S7yxOuqyIAnlgd7DoR7ra1UnDtQVx9HSDwRtQD
0+ZcHKjCTiDIdzxxQ397eAT7Y2z+HQvn3SemlJewddDte3cESrEnswzxbHNKHjTIB7R1UDCldfHU
Q9nBOpfdpxLHPEG7KrU9b8E5Y6peHV93scayGU4Qb+a3X/4Phjvdpu7hqq5twJmoMrv0cZi5we53
7MI3cKiWXmsjNMkcWQkXErob/MlaonpAYkvUR16uu6/zidBo8/el3jaQNkstzzR9TRTp0+TKmWW7
EM3c49CIHed/HqJ0g27wjlEJLHHtAfMas1HI9sbacqABIafKRuN5BT9pCDIOhDaOXMLQh9CCMCAJ
fw1EC5R9JOl6WPzrTkPz0Syzlif9a87XIraqKv1z0Xxb41eIaXZSHjfPNPSvnR0aqNS6rrt1poOq
7XEyWgyoopfPy59I2TqrtUS/Ns8/IDe0d0kXiH76e7M1FJTLvCy1ETP5ZRh7C3/Ul7ogjJS2tYv7
PaSX+sDttkuOYuuRkWV1attnj/wIIe7KFsQylMQ4FBAqBdrTpGj60WP/lM/KDDPzROb8OsnJO4ko
4I+qixNhmEBUkifl9aKFhH93FH5GAe9IAuTyOXmFLZPTpfqKROFA+tN72DMg0J2h8M+ziwZW1Jth
zgDOv1jXttsO1KS2nfvgpp9ZCtgngR/Fg6wiSZ6Gh3uBEDlMVLrML9K8fOYeL6s9/wHwXkP+Y73z
X/jJsNRjX5uLr2S7VDOoHAPHvO1leh37s1ZwmPN6Y7xdhpPN5YnTU+ngp+ovOCjR47qwf5yOfbgT
SCBTPhQIR0YuO2rEGyTy0Ntwjq/4JdtBl1P4JdZPF1qvBbaagjkJ6yvmL8f3RJKYysgq5njfmt87
HSOAbjwT0xXSpTpZB8zmsCZnWJtS/VvB9E7EbEtcdxcHck45UljQBl3+FS0tNIGwcqIKUTWFXXTB
zzmHUjS7KxgV/tsVp5vHFMZxdgmCfqiyORfwVxhjrxeJjfClMpTSz67I5Hj6TZ9D63GfjeEn4xjJ
unf3TF0PqkGmkj0csslrSSBreUNImp+30dizMwE/mJt2oaoOG7eNFTDhuIP0UewqWsYqbhsFJmXx
a6x53p006i8nmM4Ni3Lt1nmOMz3ngsrzThnjNkU5qUtX8P221YfV0Xi6tZ3GELROz5Rh61tnpgfr
djz6umn5opG2L6YBX67oPPDMWBQzG0v9sve/+D+2LScr9RKzp3uDJa45yY3ihUWls+UaU3tvaLZO
ER/dfn6+nqlhjYN1o0C1pKG51mqar2IdUDxTLqHf2vvzY77CgFiOQRKAXdIomdT8eTTYDz2MIKH8
lrcsBytrJbbDvCzdGt8eMzmkL+qep2ySH8gcmCyOOPi2b4wNsMncgUNq9UqaQkghUy28TctBUDo8
LrolkYBkHzljnKbQxTk7/x0Or2BmSoNQJEJyrwETsFlNo3fpy9Axf4sbk7CR1vaF5jtEOssz4Arf
Mp0B0Nd8vKDiUMjISbpQ1F+qaWTbP6qzRclC2stVlhpvrrBN0QvM0j78PWh9Gy/dRSSPSSWkvCss
+Zl3YOGjekSI+w4BEyYOJmiqeTDG/M0Aqb0x8j4LjakJADtBYZDu7o821uos7uKbxetOhfE41ur3
AsGEHLA2vIYj4Rh4u07K/tPSxMK3vmGxsVZe/paug1kwIrOO8avcPQM0o2yqW5HvNAnaexAVKPYv
ahZqXgIIdfrv/IjVTcu3x52NQR3xH6DZYW/6C3wIlgsBixYLpbEoObo0Dwrr+iEJr/R3b89cbGE7
qh4qIRamEAi6tsSn+2NuwbZIJecHm9XVNjmJlW/nEi+lYqdT2MlnKBwUyxVWx+K1Fodj5BStkIY5
0+7u1HC4S1uN6M0p9QUD18rOA+qdEPQBr3aiTZJrePk+6vN8ldhbAunrTEn3XYLxBhO9L2RaJu4g
5zIzp575UROqOsu8Qw3MU2Q2NIs/sXwRG4qfyAXYVH3gZsHpT6hFkqybB8GH1xRStPPtCSFADgOI
kfqvTz9xXEBLrWnhWkuFFkQ90I5eDKvPzLkvLwJehHGNJT7zdXL/AOM8Wv3UPc4nkqmlNR/WJdqf
J0vFkOpzohZh8BwgTQKtD2Sf6w7cHac97nT0zhcxEVlbTXEyk5+p5vOFQJVCMorprbCyHJ+R3uEd
xD2CEaIX5AcSPE7lP9rir0z2PFx9JtxP5uupkZMbEKEXr/ykWTaoMRwtlHF4RwlcRrJ0DVZu5C5x
i1woAiDq9S6ERfcqCi47K3Bl9xKuUnt1Ty4YVSImfFMk5OoNJig7unJ8mJl8tdkMIx7gOObbfMEc
tD7heHKTVKk8r8d+vbwjxQVFtdBysxtYy5g6Sqr2H568VmEYSCYSPBoSPz0pvOEsaeWxH078cepU
O3pi+l/S76oCuUO9D6skaKHeBLWS7k/QJewpJCNsNmJem9rbIrITWhaH1GWxbagQPIkEZPrOks6x
TafA1on8WUjcmUdyMuObmOCXjOsZ0E2CisqhHLedXpoxb3lKoAXxUsx1JwD8D5tSTgcKVwtRq37i
1KL3p8l/E1bWwL33y1lGB+XaJ4a9PdATfDtT1A4Tgg5xlf8zgKi3nqudIzUIle1GMPHNqAwy9VQy
0F7vnLl2/h63cSIpdVV3sWsbTUA6HkUFbCKsVPcns7KDfuE8NjrA1UJ4dFNxhjf7BUivjs4S58CB
/AdT10iTIofK5ijS3ygY9fhEYhnsFmcGpzlogleBRWH8nsT7JoZzozK1kmYGiJFO91tWzjiWTU9e
Rv0ICh9sHPLwN6Xyj7+CLhBz9JwRqffZtZcmxar0wky1FD5CjPUgVn29GKLiid0pXPLgFVB8AOmV
gj8beurrgFf3CyXc1q7P5yQ6eZ1CcFugBot4Sj1oXK9ljzKtLtLzGVbpS5v+bFmq29LGDvsp0NJa
VFCRH62ymN4ezYnzDXq8IM5VmQoV2oObeOoIa7GGLpCWyONuds2jKI28mvpcd+NnHYjLnK1C6cto
+vDu1bgLd+MWdT27NCSrp4yME4olRKjwXAY7Z44F08AC4CNbXjwpJ9PR9eSija04G8Zyz/aw53da
gVM8ax3GlZKoINpwFsgTmdcB64lVCPSDJyKtGIaklHr1GnHQ/G7JCUR8mwf3yKAGBYR6TkzA0tr1
4ghNbzFbKyy8IRSmChskOLDh4uIusSxAVc5CDoh5Hrc85/tVK6Qc8OZj70j9dUISkpIQRRH7yYpI
iWfqnafqA+d/ei4wbSkFEc4LoJCEf6j3w6ABP8xZxiVPmKtTyTJtcL3AYwDORNtWoTUkx/ir+p+5
eyDNcC5CDhR/oF9Lk03xIwGhTxKXYt4S7VAT5THuvlJCfYHfjGA4Ug7CI5trvo3pBGA17dVns0MS
1G7RCpAMJGzf2xJNIaNtdpH0O4cJd/vsm7FrooHmlpEsHPAO7erWmPWcm2/S+Ek2Z6/CsD2IdDjV
ioiSZR1RPtK4VdbZHOlhGao+UwxE6id23zGj40E1Vl7a+I9SZX/gq/H5fAm0fVRCNpgnLcqQfuj7
XgsPol8v2ENrdNSNGptIon+trnT+7/FqfWPY9RkFCOHkcOodbGKTBerhRQ3Umr7ftKeLyP9VRkSi
s5rV6e71CHLOReWPcTP8LYI9wPMsObkPyEAqd4b7QxOcqO//QkNtSgV6cN4ptfDdenBhIjf8FHa/
Gfw4FHkgbG28hLn08L+UtJr8gpWemUIME7rw6GjbN2/bO+hPlK4a/sm9RM+paVDQTMDEpfnvVw23
DwjOHcTIggXlqm7Iof0aqeXUxLvWso5vKon5vD/wtQ7Jy5Ao3fPZFuxI/OuVoWSwu6D6OPNdYKTd
CC+4bzHUf81zhRQ4kD7FqBYyhQUnA/d+2/COhbOt7kS0eRMGCl7784mK4DiKMo2O+QZHKQf9I/jd
KI2ZS709uRcfcBAcQNKj3RpOs/9GjD7J4vMymI2EBTWowrvN7qDLeKXNGriyu50F7CDHPR/qSsgR
/yc6ESWNWQhIwCp9yLao3LkUSmK5+5FfB24hr/lOCwksuW3JMA5xM75Eq1LN3yF0x57Dnoz02OBw
HQ9u8mNYpjpALd5ldBvW/IzA2OozcVW38v1AJ4jBIb/Dnx0kHojgUwHa7xkZtifjUv5C8OcxyyqM
GPVzVTRIlgZ4Wx8GK0kV72+8wMK7nTRDXA2A3lc3RoeWr1piBhMVWjeKuFu1C65B27IctW6ocT/T
jd8Y1eoEgZ74AzBbM4KjdFEsMyF5/Ql2asM5E6oCRFK+dmjBpnqMVyYcvHzx9BS8svipCEvO9EB1
Uu4GvfKF60o+8RhOFifdmFlOOVidy0SLHALvixlqDwWXAT96o1iNKv51kL5er3HuhhH62GciOHZ3
WGXwK8nH9qJsJked5GA/8/0ZOtqzjT0LfCibbnpP9iCEyTsxyIQ2T+UAJXzT7KI2oeaqpBo73/RK
NfquuCHhny8nNgpQpu5EwEMM4vK5WXDb3s99OedQzYUIpu1LKLruFKEi1kgu5W23SPorIqw6sabr
0FI0WtJNIqknqbNrKW1D+173N19hs32i+c/0EpHxmSNjPax2K4N8h8qVx7+S+bOCgkFPA0bXR3o/
46tQz44qofuAZ7m05rkO+m+0vh3imtPY07hu5BFYtT6X1kU8w9TDI+IyPGn6qaUrDh4aZOd8ANwH
wicj118AqMmgwKT1nYhIQFbIWZncEpL/8aIa0hYUiqgm39+10tbwg2wBMTMpPgrwoPCTGzX38l7E
t5oaX1JagcCW5SdKHbhnnEUQDIGsAxectZGWc34SYO+9Qsr7cmx40SoGvzvC2C6hnW6NNctGmS5C
UYLbvwakMw56L6d96uc/acY1vgS3eBnEHePuQLfNiz+Cd5U+IcJOsG8olk8hjLajxOY8oHCPoHvo
ZIu98MQ8Inrc9gBkbA5x6zVoll3cFV4qzXfQ8DfV379zzaL2vcTtbgrvNz6x8cya3vg4S8t1Epmz
f4a4vu2TrBj33rgtWDgArTa+TJZyE7MMkLy1F9ZLYSUs7o0HTDgfGhTsr4IGTUMlwp4sWk3FF0MX
mad3wsHHm4z+uTDTOsgVQDr3Z/cVgJi08huW6yXHLwIDqS1YxurIIWCmCKqAEdZroj6Nx7KcyAr1
sZc+Y3Ah7m6sbdzs+DZ/apEXcX1EtWpyXFkeIepW+U2At9KxVtTir0Vug2cxgX+HyMHgjCtl7mup
HHhHX8DyzaL0Dp8ntOQV5b56HE23EX3XSA+atFQbOjA7dwN8FrLskgAfnNRxeeCbi9Q0hRoliQHZ
gIJgYKmiWuh1EWPK5o7C9zjLXARpTLoudTUO9iV96++LENv4aqN8JnnCdCJTnSRaU4omT3VS1PMM
ccxolwuR4e1Q1tbS+RyfJMjfAZTfmaxtWajiVdShCH688f1NpNzM38y+B/ggvIIaDzIVNPXoGDpT
HAskRhE3cDotaVUJGL6ZPAvWMxDzbXZSVV23uziDlt1QwVJZ9yxz7VsYkdcIGVGFMEdk5G3c1UH1
yW8vaiv4I/R2ai+U2Cao3DJmJ/4NoFMkQWzYGulF0wpp96zdZVk43G+GTAkRLGTI4ObDEgyw11aC
XNG0TvYzuec6YL3rcd7pavtpXmPajKDjkei00m9ZD8Thr+GZiMf8Vc8PQ45UojN1rhCp5szmSOKH
EFxpTmrw9RyIAmQHz1r8NxwuGQ2OcY/DGmA5KDKOnY86oPJjxNyosvQUHSM+WwxCFpmeaCPg8md6
nhrZhmszw/WGswCZExN/+6muJMHE2XfYzWz6fRNXT8cW8wJatpB3tyiN7rdq2EdIGVFScul3i53f
LBEdmxdqf19cNW0ZZaOchrC3Qu7T8cKa00IUuKAJ0wq2leDWHotFfvsc07snpEz/tHpfDdL1MDhk
lAwMo6Ox4tLcLM+QhbAt5jZ2eY0xoKN/i+bfF+dOqYsEzyKqsyXmavM+ooYStUq5YzzR5cd/S5r7
tyNA04YC9SEYXHOXWZXJWbKHDhIJcwUPWHZCfBmqV6S0mUDK9TobtImBZ4f+HDCFWziM7HSAGuyV
d0XKdPQGIyreHtmw205BX8NgSPX0gOPgwdV/IvDLvNnE/90Igh+mQ7HY5QJ2zhDC+UNkyq/+dQ0I
XnU1u6abxr0tSngZbeMWl0WYNI+tqV1ppTtEnmRJLHssxKShq8cesoVk/PQkb1D0T77fOmbDavmX
RQCrrMwB146YM8BZ0oX0FcZcPExttTKcEr2IqE/mUcStteBVllPPsAcYwq/CmFgzY4lpAT6hR46H
7+z3K1wL8fMs0VQWoorckA9J0K2inFe3IzID2DF0M3lpGMg+fK94X/9pasnHj47yQCUa/VfuJmbp
cUJjbimO1Hy5SVGPMPtSETmP8RvbNLolxc+1h7uFBSuy+EMJpuK08YsiXK99uR+Horp2aAKUXb+C
1x5nEhK+pIjKCh27f5DsmTe843ImbDhmenphgnS/8SH/B5VXB9JNE67MV4KT16phoW/IXkNbv/94
LGQ+iONPyEjvMse6+HT44F9VOS4gftdhcEJLV97+Bz9JcWY5iq+IShhkyhOKe9BH64zAE07ZsZcN
fHchxq8aJtZ89kSMEF9RiGvL/f3QB5uDi1FyCzEQgvD1MdAqc6/dXdN6WxBgyJ21WRm05BK0S/fM
934hPxNMI3rLLctKWhuKCsMR3bWO6V+k1z7mZupbp0S1ch0IfaVAUnG8lGI7yL4GVekDOkSCsAAG
1s2GqFKyxgE9qMGnDM2z6hQ4T/+t47kyRIl1313JrEYWC2gt5HFkKY+x438+I3lZYpNcSotTRCtT
305nO1HKb/bqsP0IDwNcOsugDb8LRH+m5QV4biK9+XzrwSaWSSw5x8Y3lVJz3FgSjivwQjvXnnnj
/LKEpLD8mNdVmZ71qZP6YO0RVPEqcekXGXo4qiXfgddNYKKDoKeGrSV0aU6KaD1Mjge7ibJ3QeDv
8EdbnDbA+8GCMyz2r7tMEQwieKkeEYuMrFrjq86yw4Q9TykKhevdHiXuK4INRxUl5jYZs4kRWmpD
QFUP86n8v74kOfb4TTvDEwN1H/M9gP1M8bGifhH0pXsVdPndqXZhpd95o7tHK8xlZKrFgewEetyy
X6G+csnOpSttFnmR5TKKsQF00Z9qxHP0k2qzIEvbuFOMGCkWaV0MtThRIZdJIM2JhzlNzBdLRIk+
OLPbVmEE69BEcdicORez2yiWqTHQNwUVk8rZKoP4ZkxhBhEcT3/8PBbKdIIWG9NnV2i/g5vv81n5
bekLH3g23RB0KujJZS0naxgC6krdsCg/JXtLj0zzwtS0O76Z+qIiPw8wFE8WTwtf5z/SikVwiB7y
nrVzIHFz1o7QraNjd2/I4gd/NGATPnIzTXn99SDg7tw/kcNVK87I825HEix3YQ1cNv89D2m/Vgkx
4pKHR34kHLjBjWSaq5ltKfZkRyJk6ZwnJF+CPSkc48EqE9PDs6ow2l0NF1cud662dNKIi4etbTSQ
MEFEE4XBaXY8RCbwkFa36p3G1C6dCYn0JcyFi8HjnjrcNVLkziDR2qVp1ZCK8BcaH1Z8BkameWF7
D6xA3yBU3wamRPhyHCE7q+HTE2StKxKJ59/vDR9YFvKDHbPwV3wabQTYoZJsgkS01HqvXgRyrvbP
TS++lRN+ODDV+Y0Lr06Kc1PKN624oNRtMN2xFzVdb8vqdyM4lfQVeapfAmtO8feW4Oyqidu8Y0id
2AQLNmw6B6Wc8KLuPqVxnFTm9oxotGDMjXiJG72QjoM3mzz1XFF0dwxxRVsYQan2BImwsLjUrjbk
bmdMtiUHCxBH7Eu3xHf7QlZ5w1fbR/2i009Pz4rNG+JY8pi6rhMOfNIyOBeCn7lEj376b8Qp9hYT
R0ux4+6emFY+QSdYALE8Cna4Ur9wDLWMlCGaBzU346VP3iFYk7+BnVL50JtacxBsuTK/KKVMFIlo
znwdyu4MspjmtcADgWu4leM663np4ywf4atBWAgHTAEMKl1e6C8KyYx+Myk6QXu0DNmL0yeRb0wa
tUljcZ4MBbbE1cSQca0kUEPEXRbJJ8S3WELoxMaLzwloqqulTdCA4Z29dBxH3fLHxtQ6CDFr9IiK
2+X4nXnqf6aZHa0jWumJ9VHImpfmEaRJ02qdmXqX+tVD0jk1idoU9x9fR3tEZn6x7+sv0s38dmKC
iGtDxov/JUZqX5d8KmTlhTXU2TjrBzthKTs+zeIfZj0Gk1q7KcFVAlIOQq9rTqzURB7OBT8TWPNk
oHs+GwaXDhiE07CxijsSvcL/d5o693JzEfVyLQ+2gmmE5H7UjHcJT8ibLBgNc/FuSzmWNNzaKVFy
gBZzqmM9YCO4HDSPbosduh4aox15+RR3lLaNnj7DYkTPzriT3v82hDV3D57jAfuRfULmrBERpPZo
YNYMwjLGQQbUgw6W2ixeArvCUeTLNfmcKUv2faqhQwZV1le+xHc3le1TjMil8zb1PbrB0IcUFltY
Jp35ktpxjK/YGIcODdoQli9Y46Vk7S69VEvesp8P6X27T5XihRp23WkhdYT/qzxGEl+I3Z56IQJo
4vX//TghpdNrTHb/M3BdYGAd5xfv17pC7xMTO4g6vW5bJXSVAE54TONwzl0Yk/a7Getg2kJ5Mj/R
6ZzMvQOWAdodNW41/2zGUiKM8qp+j2peILiI64TaFEYcar9M2pn+RVTNPMYFb5scI8AtG2gbzxOY
lxhv/t176ivIXJ9fvemRHGX96dCdJc9M3D2tsM0r20lqVe+0CjcZxANVtweCLfb69znY2DBsCCLY
uEgxMrklCV463jUMF5Bk3Mq6W4opRIxIO7x05tPZ4VaauOX3pqTvf7fCDBz4KsFh6GzTqvA4SZDp
w929HDht4LLmvIKZ/9ZBPegXU6dwxQNn7j0PoNsU/RVgzXfOGkBmEGL2rYBVw7VCK0ZC5BJtm5f/
11+uvdtxek4FAGXr+Y4XPBnEMKJoRc1WuxI1q+TUlB4Vsn0z8OzXPwJWJmZVgZpCSkFD2DXt9DpV
RwUj1HWoBYKSUOB7W1iLuuJOlFk46ZtWrg/Zrkb2COmYaBkBcBnGZxSV3q2s3lvLIM4QYtLACIdq
rbEP+8j0AvpDg5vzp5l4mEEteHrzLGSLKDrQi8Fa64f/GbkCagZmGOnYEKhOM7fuo0sUMTYCl6XS
uRUHiNcrKAZmNOKTB8fL2Zl+tdF+mR0um9YvAXuGIW1O7Td1FkKpdsZe/6cnWbSTUmRkS+832Hqy
GRi0d2TtYkt4MCrWX8NJXn+/Dx+E3LcRZxbD/xC8GycnJZAOSP7XRhIZWUfsfxSeE2xEHbUcES+U
XqCCrxZ4NV3lnAey5Qvymmau50StZGtzgqOlg/tdJD/ZgfckV04Vn61xLj/z0X96nmH1GXdWwssU
524s5e4icXWMQ4V6vycltv49461nGtKu3D1wyIb+YrjmRhLn3bNNT6T2mNbpXzDrSapxC07Cty/0
y5HRHvzxfNmfVAOsQu2sYL4UuyNI0VyGue9ru8i9ZZVsvnmfrbF1IJQPDc7x0Ndngz3KkNMaXJfK
J1cg6bHF0+a7GDCdvufINLc/0UHFchE7AuBgVAAI/m1UvcRgzBp/j7BPky4Z7vG/RZ917y6j4PfW
8ScFjv0fcGrZhOq/WD9K1SKs3ja4Cwo7rLaUk7/rM8p2ArYoxL1D4BhN8xeEphFOGJ7ZrXSO/E5C
kZqJURSXiglLfyGh9R3c80xGQIqbT69tE0lqzDzMuu0Tojl36GtxfJQUfCfNQG3AZ99mb09xo4dA
k4DYM1YwtnAOZqx/zh6eUWkBu/BTSZi2TC36ezbjdwCS39VySXdgAIsRZ6scLPYRbCsI7TaQMCIT
k/zZ6w2FLjKtZVibOC+VrxgABKzDr1tDfxWpcQTQw3mdSHfSwrkhd5Guc067VOsgHAAx3SSx5ELC
EiKlZZVSrKm30W/UjVdvNPgh1t708aUoOznrSsghc77AfQRpA7SfvuxPXXO5Q/EVR2l8A6EBQni2
BQA17F4KuNP+rgFVwesG10G2HHJ+Q0kilmhKoruAxpmiNlCZ+doJMQ/RMU9JTIq/GWj7aPGUHBEB
nGBsjEYc94J9gWrdjtFekUqMpBYGMqoMky1coBF7zOlO9oytVzDbPttLrAY+0gDveJnypHOqz+cQ
K58K5Zd1bGboErLMzBGvP3iIzi/lvXEyQQ7B4Qa03u8F//Ntzk9r/7+GstBqEF0q4z2e/XpWObd/
dtR9ccN5/NVNBwUGpj8UBuNW/wC4zZOCJIMbc5ALdU+4s5N/H8bmPZ2jsUXHM4vMr04gY8+/Yc6U
f9TOl3U+yIUVLwDEaNyowOEn/j6Xxp3OO9etK0tSJSnaAJV1UtlT4r9Uq/1ZgBa5UmWliecy6x/n
mTP1EOt9wEq40Wiptq1t2jHkDOR2BvzMB7jJ26wCFp/N0/+YkiuiZWsVZXtuB5EkWXyVgMXFMUg3
KEB8p5o5gJVKimoQWBix81jqzjk/dS3kPwslF7VDQAdE5MgNRVWKxrdF2MmySlsNbuxUqxn1AOvj
VoTqfdVFvffnFJaQIH1Za1XjZbt58YuKL569Z5MATBEyvT4xew4uXQQq0VzvmLgLRkal9n4PrgOa
OHiwAOQv5aTrIbHpLEr3eo5lDO98x9qNfkgpAzU9+RBg3tvqV4NBqBvL2nd7dDpulczZdQilrg9V
H+n4GHDfoMUvmK+SV4TOZyJV1tDqECxR706tAIv5JEosY2PJcaXi1I/eahFBKKVGhSxEg6M6HwGA
MzDprJXNfXpMRurrWLjh9V7EJzziYhVwId5dtI4hEVzB8VMLAxYXkkSO+3QnBz/EFQXlm0qfPu2r
spfjkXOMYH+0HL4A39BfNoueJxvoZ9/fQTumInkct9XWKoXqGtAIL0Nmw8Xw6LSJkF5zzGDlkRim
9MpYbjZu7wqeGx3fQrG4FGXMjeEwbGe/cwGzX1qaZJoVe6Gg7RrLk6mBm6HochoipYI6VTqDsM5d
f8MNcqJK7NQTyy5P8e+KQcsZO7SecmFNK59/V21oPJ1jnjjQmml3s3oc/sAYTST3i5f+iJ9RSBkW
SghF+nRhJmswGDreZwL56I+uCB+CXuvCjiQfI6/LRIi+b3ZwQpNJV5QJTq2D9igfooUkyG/A7gd7
C8O9cHssISmBy4mrNzl+xZ6wnEDDAmHnpxlpmARqefmhPxGRToBLnOnpO+mzUNQ2o/EdowkJwP6B
50Nb+yPrENEMy9mqjqO/7tELkEstxxp4xn8wMkISHqXgvLQ9/Lj7SqDGTgSPdf9APwcmLA2QabEK
ESzPpdfe32XFSwTetZp3flVxUjk5AYuPytS+k3JcQxbgGWDYCioQ1jd1B6YssOgt6J7O20JDpI/y
fajVntvdxap42y/8lwz8NxfuyBS5trVoF/Z1z0tLciNg6uTmJV3+ypuBnQkgEffahYgf/Tu8St6B
246jifaZLLeNeG/ZjT1zPRDB7zPuwiR9x0ojwgsV2BO8HKS2YZKQ792YFG5SLJE2JLVejcT7erMn
Rfvvay+M4d7G3FAG9SB0RuW9YXqrmzcwJhBUEvAF4kU/rUmAD1pwYHfU4PM4lYv1x/pbGcyR01RV
LRnDBhjTh+wW+UEuKFegvKLMc9QBY86t/NPl80JliWnPkUTxffKR0nABFpGOq5Rn492rWposWf+f
49HKvRdxq673jVDff+2gDNGU0B+Ou/uuleea+jGo57OBcs4FMmzNymZxOzq18mOCks+xhKrCnHVS
etzRJsJPiGW8JVdL9IK68YoscEZ6coZDD9C5Gfan/QqdTamL3ON93OLF7Vm2ch0l09AVhG7yTVU+
lEw58DLhj1APOzMHESDlWUtJxGnxiIAbTKxt4jHrZo59VCCGQwOOrxhv4BxLsRErtYoIhmdvp1aC
oRZO7GlXKk7CA+Hpub3gxsx6cxd51Fp/yciy5M2vdB4pxWNZPHyjJ3vjTgJFjdn2odc10WweHwZH
PW5mS8YvzNWhON0XP1Nb5RHvvNyyTViOMQlOYOTgVbVmMc+abcdQArrM/PdcXxdF3ANWE37vK+OQ
xR69B5Cw+xk1GvDqmsYNU6Y+/SLZ3ViH8bhjCpf9M1FayawMZF3YmR4X7aaScVWpqehDcLRSUPSk
Zp7mF4e+jIa/nGQbB4jueVAMH5rm414vNx5Ru0sbRDEhiKu7izuy/sjUqldgptRUi7rz2EDB8ncG
/WyIPJAJXpRhHMbyh2KfBmc3noOrrPM/zRXr4rFemlTXS0P+LfAeo9wlSYn5y8ynQnhz4GlZsCd+
bf1WpFvPftetp3K6kJT/ttL+Hv3yJY5x/nbtN1/Q8e5sONaXwgWn9I/M3rzvYKQtECBWyfb+7id2
t18YDcbYbS3Mog2ob31DL+QApoe4u3b1BKD6p9tXD9hEcmDKQewE+xrS6+NEYipeSr09TCGIVwM/
DAq+dPLFaqiOlTc0ghawlkqXjDQ6QTGiQ38UwOi8WOfLWS8yX4o52tG2oEwPu0aiVag4DYRV4Gro
xxk3b08yhpIv1/FcndPxqtdHYp3S/llmwwHyZdTWd1KDR/n0DIMDyo5jq/uf7Orh9bciegrRsr/R
UXZd//ol4JoUkLIAEdSyN4jTZ1FnqySbfLztv8fJnX8OI4R8yWv5smdyewcZ0e65uczLNJhF8K9H
oQdQ7pkH1x5Ho7aT/42gBpPNLs2rlYEgGun2hpjvb9rGQ06chjpQ0pECBm67IY3ZTEQd584dns6S
BciVmkpu/EvUUH6WCL6inZZclM4XqglQCB3m4nzeqBTNsz0wicejPiMbf55dkkImtp5IrPlZk9o1
FLvSz1wi6jwWXIf54+tYx8S2rFoWF5vjAT9LTmhRq4/zZ9AgsT76chOrc8nYvvWIA6667WGx48iL
v8/WyeHnc//26AOx02DtrWdCkPozv5KmmkkdmAOjxDuIesiLqY2RBsFKtDhbDSzrBgHtSvmQ0MpI
nI0eY9VuTT/OKb/C/j7vk+IXsjJOJItBCBAcZAA3xpqgzcliPtxqhFXfU5HY7LYm5oRG5XIbfLQl
Nq1yLUSQeqyoMUN8q0R7XvJycyo8E6HWeyQsvmxMtiTmNqAvn1tg1g/Npb5gFsQznqdmTbZnPksQ
r9Vt8yXmgFyVEIhKW/77ZKWSYjnZKbxcJ9Cs152YD1m09xVUsMcDJNK4+aMnuHwOskYT7EU6y/fv
SluHOczKjc6BHWG81slcmqOIdUf9IfbeyLcHXBNunmcfFS8g2m/DkAQplz141GkdC9Joev9us7QO
/YIaHOA7qrvAH87QWel1Fqhmdm7OxflbTLhJZCrCJZ9TqJkAnV3TuKvSx4U24PMHYka7s1B6qR1B
6MaU6rrFLkGam/xk/zu2xVOcqI9za8KNqq+Y6mWcwrtTyYBkf64pjBPu3O/Ws9rphqQk+dr6X6HN
I5xpNiJtgpBafSMcFEMkMQIM4iS12WQgXLKwCzj/+rZwabmYvA9gL5LGhuF7qbADDGDRdMDEetGj
EoyIYO5gKNCUgK/B3oicFfHdk6onmi6WeMdaulHJPRz7Gj9Njyp7c0b02SfsWtdzcrJGcTixJgoK
386BiMFxA0vj5zrzsskpVntGVoPW0vCvMhKg1QVPiMzFa/TuZdv/QBqC8O83kSf68bQO/oG4CkXQ
TzKbU/PvFgw3BaqTDhn9UyVd6gpSTLOTt26cdvFi4o6Xrc++xrRf1A09Dp4AB1vvjM+YGg3vUBBr
798pcL99NMOt4BeBzddzMkOA1hEbi1Z0nhNd2rPIkI4Dsa2+90/jy8X+OsphWJtsrrsjIffWVTCN
lfuJ83LVGJfwtPmT5D343kubYUC2Jq+KdpZlgEWbhmc7bswoJj2/tu6XXz4CDdb/k2qkGDAkO/nD
2+HHd+kY56aT8nL7rEtaRpywAFMMvhkBD6xIaxweQzVf+Sr66+o266yDFWV8tH4YEFhiyR+D8nBU
CTdUd77s+wcfyU26XhKJzagmdZWOQ13/Uh0wfvnrs1kaw5wPxAmEq9/mucaiRTwC/3ybn6m5wjDW
4wJfooxH3KvWixMSbi/5Dg2OOm7mXkDRHhxsfW1GPtaWfefl5f/gKxTrnhNd08pa0mvOUqaq+Arm
lLGUMankri5BvuAMzGpOQOsoHnmtfDSqRkkhRT6C2fdGvYZtF5PjbMgcwQVuhXHbBIOX1+8sYMvJ
X0HNwXimaBq+QgDMj4wys3jVn2YmsR5Z8tE0EaX4tzWS3ggBklqcDDOxIrGn6rQb5SzDEAqHsRbw
N73SotDhUJntyau395t6UJHVNwgcgiUX37RqP4zxdsFSvgATIreygemrtwUs2ePGqDzCJ49Q8ckr
s7tATr43PJsSu9EsBdm3W+q7TmTE0wYG+xNuF8nWzr+SJXsBFsT5oiAqGO3FGJcxSiCUdvXO3hFe
pajJAzQceyBhvIX/bCqsjf+w3roRUWzZolRoLVxpCFEmGw1D3JCUSr49V8VSJels38a98zwWe3nl
ukIEZUm57+5/HSIOp4Kq7AgKHkkB4h3otZpLz4OKOeMq1xJwyYivuOBfyx+Ywx8TO3OYmBrMaxsy
yy8GJW1QruYJbsGLl/zLMrq4SDppX04XK3tSJSCUEHtZk8b6T8poq1dQzmry4Ukue6k4Z0h6MLde
Kl6oArqsw0M+KqlAk2WmTN5cTB7PXahT0vkNTVsZV7zNOJOJmffQyBS7Ii/KDWvX12ZYt1NDlsx3
WiO8fZRwGEpCw+skHJPPOEV9eMu1/ghsgZjcP02Z4iCfOI8w+Dn46jPThIoe4KKVOD0WvY7S1tPZ
L0YJVuBgT7CC/QXSz91OZEkzrJ9Q6FiZIurrTTLoBLj+MmM+t83esTRurNLDgrPJ7i9H59RH2ScP
z7qgBKO+Yv8llFHgr2/L6JatwsIKBb7F4zVIH8lMikUofckeZDM3+YEKDSa3mKi14hybCXhinfxC
8Fj6W/oP47FcbPutM9QoUX+I7yQkrYJCkKkgcEETnO2im6Wbgpz7RYjDKRVnJNjK7NSlEaNzHA3X
Veq6zlT+mEHmsVivrJsQ++k7eIsdQC8e6y3T19IPYbMdBLMgfs06+N8gjxjFnEdppLX70ULRfyk6
39pubR7wPJcbR5fNb9Mj71B9jQkSq9AjThfUw9xLWrW6K1srhZwY7Har+TRu+9qvi/iQUrl34c7o
5brlQU85mNCLeCP70mIAKrTjU5bCIMWN4W7zHcE/KLYEuPJzV04AVvizii3cw/1U5SO+zvpyuv0o
pSk/eWxoNJwsx3elNXcu3otdvJIFSbkBlUAZYwxiZBwVdkWHDmDUVhGDF8GUp88kPPIVzMMwAYZt
dIY3/fYI5fnMUGsedh/ivit0L9j1i2rHDChmdxfy3oUlYqXPh5ABJb7M4W3nFFzWrG+UJU8F5IMN
po6UYz2Ru4qkQOIvk2siRGxCk9kzblGzl1kHscXvsLbb7LHXqDD4nK/PlK+cFxeji7CveR4obD42
T+bwUdBMK2W0lYTFsd/zM7BXsYmoOGzAKKeL44YCH7F4twSCW9zl/NnlrR2L5xCYnmciuMtiQ0es
DzzrAQpb4Pk8yubxUFC0/XwrzWiXhDCofZ2hz1a/kLTdu6WUHLiVJlPmil+uFsMUz6+0R1aOIwDb
OtiaWs5VYnnzB4azmfFciXH/vEIQqIch3hH9Hyqn36XuONAQJ+uwkRZ/LXP4RY3BbsENFu+dDEzF
6lBQvG8QNi2GWA1A7jZBP5VWfNb56WFd87pCKvzPealeDnioqfy9qbtBpBj/igI52rUGGYu0Oin4
ZvG2167fX6ATas87HUau3UlRebVubH3qaeX5WpJ7b5URaRMHYgzCO9IQ5QApsyiqA0bzL6qgwR3W
OSGLBvD7iHG32pz9PQOJ5H2Msd7GnnWXRWUk6WtCjEX9lGSIJCLv5SO59+O9W2We4JEr+NP5/Mwg
+aOhQ/0VyawjAe3YHVKNR786ArDE3yB4dJ8If7WGmHwkrlTDDnmwn3pf5nr9SFmO+Ntqc18o2Jsv
BiyNIvOg+ukM6EIU6UjoPuO1tdcpCIRpDMQ91077SIn106VV0YYTU0p+oW0LbAO3fsN2tcHvw97q
AHl+RRjKw+UMO1dQ4Pbb5osiURtJjFi0ER6dzKjdBIIluQ3YgYqq/Z5SIEpIg1u9ey//XW8omh12
11EseY73f7kW1sQBc0jdMO8Cv2chVGZOUkL+P7X+sQI2QnOnIGgcX5Pxfp6FCqBe69RkW0bMwzTn
hFkAbewlRgKXIMnFG7USedkxsJX4tnraVRvfjyOGID5nM24zBAW6BdWekzvttQcITJTG7T4R4xsL
I+ziAtlba9nuA3YdeOEZV95evfY7zeSBC6LDkWhZc0OkLJUn+P4qigyC08K1mIhxe6YKFU2MKoEj
DK1C0BHoEJBdqcUKMOpjWq6i02uRqOxxHgvwAprlVeoMgXzLSMmOTJ35UdLZ5hDtCM3vWLLkHxd8
U9DpIFsP2PurNg6MVjK+NPbwbBR2u2KCu0U//wYNSXtWlWHTPtYdfdRvc9dmmhLFWw4dTh/e505X
I+7XUXJHWk/H88TZfhKLlBV1pNbIAY1yAIkZkaIGiAQT+C9hgR/776kz+m/c40b5acpHXraEeH/2
cKAl9MLUVKFCh7Cxw7Q880T9MgY880hXfMGTd2t8KKlG4yIz/ex+iTd57aoNgZhI6/9W78681BH/
JknM0QmwGAsHL7NtO8wSolOihnPUcJ719QtkNZzyVvlgpb0jlR/PSYGRRdQiLrIag/WQBoyjW2E3
EPEsOFrFBaOmZiipa6LbDRDKRxuzZQU91De4qGLS3dc0+uIpllrYvnKARCP+rRgIvnYM6KUhKG+E
76NHKifY0I8d6McLayOItNLM9m+78yAkK2fEsIQG5ImkOed6oZAd1s0lwa/D+0XgZuM3FjvNTAT/
yojB25EsY6zBTTCKYfzYN67oXx6kBCX6uFV8JZyh89AP/93ekP4zZSSpeD8qjIBHSzb2dBkNPNap
t2F+kizmM926eg7LNqdn3T4Y4IhUsF/cDY/sqcp/gU6HRi/qObSZyg3udAJ/YgVN+FjsWGt5TN3u
VXffF7vgzEtfp8fVTJ2ChsoJEBF2/4tEM3cveJveQHYiAlko3YTjaSxwZiybIXw1wpS2T4Kcyu6a
tT2w7IqwlpIIZEsR5zmQ9YQD/B9iATl6ufFgg4Iwvn7Jb4NDIMQKLKqwk6DSkgt03mXzvrpljKu+
vHDDNIYk051qDGNU8Zv8KLREM/6Oua0I+uqTyS3vcKMp4pdzCURPmVpcys5rKUVj0T29PTbBFxRT
ID4+RtWxbg4k75YTQ52slkf//O0+h2oanU2+6H/oeb9PxHEbuMRFZkc80dWvVxlvQzy7g8OZ/05n
cF3xtH8hC9tu16GoanWfN9tJQqbKTrou7sjiUUGrCDstTdR13mmVNx0YO+jEAzxvIQ1IsotECeRV
MlmPxv1rrm9VxAGGyLLMPs3EkdzrDBXsfb4xHRTs4Pb6oea4FSJ8xe2Uo45lhiOJ6k8VYbIpk3sK
Kmx5d9j9hvxuyxz58jfx4eR/4/RAAiC8/inJjjYbXWBHp0iOnxYaE3geemuGsQAjHwnNye6uP/u4
GiQhLoyAvVgWUkQxJC/B2R76Zr6awLXal3KDBTEe6ohHroF5TkksNa1Le+aLxjnon0+CmmYte5Ul
HbT7bytVB/zbJJms1xmEa915f1i/kXcDWx1Vck9zDjuUcDfLmb8FZTlu5yBV6XTZsWeSSNWUKUf5
4xqwMrTdC5svlpwf2dN4BpvzJTt7DkojRBmrpsfMjO+7+dpsEf0t6/UVdgXPdh5a11Tr241XuW/s
iABCmts5HR97jcSSMVgg2RfVo3ZupoKkgSm6SOr7IJ2PWtfQtnahL/0Sw10G1qbj/BFbytyFVhRM
LWAPlxFl9eWiN++MurkFZwOCcc7torLVvOz7DCCsf/enCW/DRAEcgw/u1OUfOeHXbIJEJtRz4Xz6
SLGvGIVXag+r4V2JdGEphnQrf8BmuDE85/g4lA1TKv0n3GZ03ISdTVY5FU4WTTnlCju9KDOy4QXA
YhSQggcS7PqFqBZS36D0mYRWXaH0h6FGvKqJ08O/p8ndnfyB8N550ddDZLwWKDb9DR5n3LmHUD7f
lZD/af6vacVdyuu1e4EMTc1S8qGrIufnlfTHtLKXQEYYSlOu7YTu9oD9QcMCyr/u/ivvlJvPi8dS
J6qFJvTz2gVZ5iLNeRbpW8XYYM7JwmMPi0yhKtBAIH3Eb4CsLXbMd1WhcRlphf242oE+6tnblbbH
I66Rxxt9v/t48uvjPGthAFtHNeef3U27yGwmFopVcq+QdxldN8F2WUlgZHF7w0pBIdeHpOTu72vt
Ji/mNUw9wS9NMW0Kf2W01LU=
`pragma protect end_protected

