`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OTe8G04mf+nOV06lOtsZs3wjaK4Y7dL+SIY76z2H2nm4GSNskmVPn+EOZ4RKL4/et25dbn9t2t1k
LNZJaokUxI0/exIwNZiGGSPfxzoWuPnlCEuVTcHeWoRrEAM4ZJzApbhTKNsevF/SB4Iiu7//Zcg5
0nDZccjPNqW+ccykQvp9qeGtT/jOkXpCXhGOVJt8sBnj7Dg6t3aE3QGWn1Vqdv0w8zAz+6KVDe9+
qfu33dtDziCx63YNkYYj5QCPzHUXhPLAMxrTDPPSN5UszjvPVu9O2iJLHPKzSvH6YY57V3V7fseI
G6Af6jbB/eCUhr065e/7i8jyb7goGo8u5ilEoA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
dFCemdQ6i8U0af0RFG2V2MCDU9F7H2XdFGNFbSzqn51tl7/yqgRA7W9MMHYK9VnV86bCpcGQ4WxU
7eMnBcjK4lGd2AkNCRQHBX4qGH+bIPKsZvu+VJq6qPUo97eE0QVsLAndHusMbht5U64C1i3lHqlK
IOFbhX6QObFlmk+/5WIwAxKmJht/ngKb0iNWdIsU3aw4OEP4RXLsb5N8zBwxcLZoIQPlQJuhbubJ
IngoK2R6AUANuSLFRt6HhegArbdnYa4vhX3wnkvQHMELTfxnQ1jUQS5y0QW2vxMvIzKqxkVim0CK
7LLARpI0mRWMzuahX/xXMG071vzQLPQSIkbryAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
mMKTrYno6wZdvYXV7H3bDEU/gschTWhBvrWJ+iaCSDHTtAplCZNFzbrygb9peTC9b2g7sdIuPcwB
qhV++YNJ3w==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LTlkrm88IihZpqptBmpaVGBOrInOJ0pAfSP38B5kJZgnHIFZduEg9ZvVV9y2BlOiFhxVSG0ZxzS0
NRZBwRmUdcAAzIMFc6llaERAn3Pp24T6kXegwCh+Ge6TmWOL4X5lbO7cyrszVG5FKdEIknwaq9UB
jwmanFid1O5NM9YaIUy50ZzyAehLglZhbZAwDhZhdTR/Of/2Mp5EIADJxaYaDl/l3Rz4Tei1OyNe
fGltZh62uk8YKtZO5Ou9Rrwt5Wn5BAya2uCClcY2h3DSTrp2IWMQOls3nKHUo/Gztzq/CknHyS+L
eQPWaaXVH+R/o+El6rcNGeGalE6SzvHGn+gaEg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
oqlSeuwoIKUxH0qpBjHjzEoUabFs6GjH2kM64g5IlZQ09rXxnL4vRI/U34GzxnX2jHjlu6e5vo94
pMmNML9aw73c6ZMJnYFDqgJW9dfDfZ2A0ZbF2u7sobpLkZMJWPufpquHCoM1eW7/trHn6TWfk1qd
RyHJu9ewoCtRkdFJ2i6vGF3brTDKuWcX/Ar1a6AlnIvDzMAo3TJdMkCadJFcrdnQ+Hh7gWrqfjCP
fXmCXby5DLoTfublvwwhPkWF0kaBSAYkJFQdIttZ9X64oLE5Z7RNawbKh0un4GEHG2mxJFLpkyk1
6A78Uj21I+xFpyZF8/oVD2R4w1dSoQOPrB7rHA==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
J+4WNvridqn8D4chgXE2AI97cxN6ZuZ5x+FoBiKxseaZ40HxWbRk9yPzS3BK98t5xGAhTxPLvFFf
v0kLDl32XZSh7pk7ABoU45dYiPsxnCht5xtwKfMXfRFgfYt9DyJkTfvyIM8yLcD6aWatjbfMJuAa
nhmU+T/OiI0UPoF6BYQ=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VV/F99bKTG+kiQR1/ucuF+cIBt4nC1urNU/Nj/fKIiQX1sfjZaJwitqA0NpWiUItGsxkwgUKpzoB
VS38qNicn22wuTSCZ6Bj+jjVMitvPVo4b7umlW43/p4bqJXVIJ5YO4nirA/bBHvPtCTSk0qH8lQP
N/ZBk7FJYItvachglIhiLs34mM4GH7eQUzZfaqllRCnak0x6SMYvQMV6I4g5ApDmk0IcE7FsK2Cs
jXXFgszU0bhAcE03xdxEtJYntiprm4d+iCi1xPpqQwb0K0MjO4ypjjEl6YOW6FQjBmGPaQd2pZ0L
3X3Qb+gT9PsLNbFXPF/6dcKsmBSa8apYn0dEQA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
DVarMflnLT9uLUFuISChhVOmE1VS6ZSDdTFmx6xMEWTS+EDibljTkCh6E+N+kzgLL+x0VFVRpdSs
sJkdf1Xc8lGKcxNkqZHyFduXtancnYc5iblHqUPdoFibG0QkfXl1xRz6E4PnNF19t9srEjtuJFvT
uxZiG6rgeXbK8mlaFhd6QQAlLhKnqP7zrzvU3ElUr8mVFCFRGhSHtcDbR0xAZDP5FpvWFTalxmvQ
3fq/sJgztJ/V6LCvY4P5cXuiBP/cMP0Qf5zQywAlI1yIY+i46HkB6LGS1yxe1TJKP95NPlqblCWQ
D+psbAuGew/MjErbHiSMIxhRIEZxqHdPtllfWA==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PzUTUOboeO5OEngHu2oP7X2BGJWPNhysL9n0witwvHu/13kg52BbuBj64UuxpNK3ekJR5lGrWZfI
7RoddoPDyjk7Ga4B2K8ZKOtQ1iraQCwsMf8Qaa5nV7dh0/3KUQEq94CfFwCnkgORXkqJJ/nDFKtj
YL1m5noyX0qe65L9BnU=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XtSuNDvM4xPUDevgmE9TM8PN+j8D1MGIu8j4dyJgVcWGmS4caNrCQTSQiXv6nWJmXuGFSA2jmiab
/NTdn2kSdRZ/55pEXqKsFp9y4WXf/R8qZVyjwmvjaLf9ANDEI/xMqEBEbBwaP002Y8+duFRNH228
eqcnjPWhwTivAecJ5QhYZSno33E0zksPljlMAPVO/SipR/zDrx4PmWAYeJh3/cYK0xvHYlF4uhpO
lcBsjqxa11w4+ylzQHPLTD0ZXev45pdKuj3cgCOoYRMWehnHAypuaOsouqZmJwH3CHYc+6vOjY/W
gXhrKyfMcXtQ1aPQH749DxR8ERIORscj3Q3p9A==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25664)
`pragma protect data_block
JnoQxzfK6c7f1ADiD9A8ucSWpkgrV9ZnJAgDdSeKVLM/usVzDlBOhF2Aj7M64+X/AiJ9p8WQjERA
GLVn1yGUqpfqYqtHhLt3Q1Olfe1tqOB1y92Sxkq9gjCcCgOuWA5nto61RTHcdPpDe3tDKxENVz4w
sThMn42gTnxtc3JZTbaYJxCWppebxbe5Jq6EOFwGUAD4IopXi/aM8Y0ZcfaAZG6jIV5vdG1MRHS2
wgE/7+XykuMHlZ8w42VDKw9vhrZeRwYAxAhyN4vCFpSZwVd38qWQZ/ni/BnqelVgfaCqEDGNdsqp
NlB4ILEn3ZxWDA8mar5/BUiTrW8MRyUO+wTcgvmv/Ubq5BOqdFecYQehZfgsORxTmmVGDPYaDr4C
nlVNcqvmf3VG6FSXtyftfo38AQFCzqZQcN7Je6VxwLWBN2ZcOSNbmrCr7SBszuTIcyz5R+aZaB+C
5yZev6yBJvcTXeB1YEFxHDAmLKpuBFlVc4xo9W9VKjzzOQmM3598WkQXHsffq6N/CWwZLiIJj2dB
MnX98u84rKlLJVMopgFcPTyhG8gM9fOCF4os7guISMS32jbl1VFN7RAUkd8SQnl3lySnbDnSZU3y
ydrS0c3NQepef88YOd91vO7jPDV2C0zxB0TUzi0yomyG0EzmNInfnalyQcV9qtVY40BKSfMeJb6G
UPaIJmZM1UmWh3+QpKyOuE6nuXbvmk/d6NFNIrq3RxEjZa3VVR/3CNmNX3YYXPLDnIN21yKKZUrS
8n5ysfs7kEeVr7zmtWtQnleglSaBjqV/OQCYx4lG+OxMERdYOePybgAnNfP5aL9o1t+adwQPriVu
GlZOa5Jel3dEfZdBONrJP9xCMjY+PPUoxAZojRSI3W7FitbtVH+WmeKnvw4aODSW/CDnF14ynkh4
vGQGHJKlh4fe48t6lqRSutI29WgBxN6ZFrgJ+J63pJuTewlU2WSuIyb9FcbKwx/owlwtu9qvc+Ds
daEMQMPs5/O88AXCaPNP1qDvQSohEtOPkfuDaSPNUT/v/xLh6XGwr9qFMosau7rZyRFAL35XZFdP
B3vnhk80CXksqA92nbFO8wUYk36EbYvvAM83e9uojcqSSntlwAcsAbinLPejYa73HFoQsCelc3HP
CMk/DK2uQTDcRNCOL11wnaVFdFuYUNGiuFU3C2VDvXR3oFcO0PrBlbv3amrQdGrxsRrT85frfCx+
pKWtjXOyXLHSIbV8ljH78jhmjO2rf/oUoqHM9Q/0yeHWUic5zqXMDf8GuzmxQ0La4Eg3yu9SdRI/
8vog7EUum46b5piyfmfw0JZ532WIev9pEgjmlZLczkXVYw27daNo7fMT9fM+wvQVg+JFWDz1NLUi
J2e6LJNd4ozBVrCJT8BF++31tq27d9A/M1i+U5DktScSmtD1ecFQD3bKeYZBc3QFYK93o0mRG+vC
1A/VG99QJFhS7+aCyGnuc22MAglv5dENdDsvZdSpo7xzjDWU3TeRjEc+UXk7Ahx2JM86AOVSrSY3
8Cvnf6j8XwOLmR9bjV+q+LvThQR5fcefe/3xUcvyvvfcP3L+I6KFKu9eRHHz9aVg3sH30hIKTuvE
gsg2NZt6ZeJTn8GpYPoztZkTaa+KgRmD1gHbQXHFGMTy95O7fCl/3/ryFPmPWRrs4YFhHiF1g1TM
Wjh1jHWVgbUaASXVnNKhyZagMuyLb/6mD1ew94d0PsoMz0ZYffDLLX/gJsfzcwDK4UufrQbcmhsX
rZWMZTO6zq+UOMM6fseZmEeIaf4XByQ7xEzQXsbjkCNdoH06ERBSF/Eke9aYna5qbFz8C7LhR2cD
DRYqitGi13ff49ZGnExGx+7U4PwcSCW8NwOc0V+m9Mr1Mn54ajLOY9kdd/DiHiQeSpHU8w4rFjgo
95NqZITb/LwvgmCezKId5K1/c41PvQ6Lotbi2imu7D01rznhh95+0z1pzHPJ0oTuCfhfSf40M5fq
NGVheDkg5b76KEUu2KitjBmHpa2NhjxwGrl0+Ke6NGaPylBDoR7VD/NPQ0lv8ViKN4doDmsllMeb
n1SW/SSKAgEfodSUFeJ6VbILBW2wyYyoVrPFEbjaBm/L9dih1X7PtS8KvgCspemM6QZ/721iUO8T
3j3gubJa6yX6TTwpAyDhlhEDf4NqO/WZmETwICFCmd2uk+Jkbg6+uA9Cj9amyZySO8R1nWw7gXtu
+bnQlteqOYjYNdi5O2izOH4KVXXZdMHeIwOrv8GdgXMDcXEvQi5gq1B7XV7shw7fZ/4Mx6MW2jw7
qqWAcUStkwm0ecQ7WC1GFM+ogTfiUo+Tx0JDbgh4TFZD4sO3vJLIWZHU5BVNv/Nq2jM/AZL+J247
GEqqNX3R3fZxMv1Jt4dzQr8o2Oc5oo9GPEBkq89LikDwQif7klHjuQBXIt5e3akSormY2gVksuBl
WBo1yKTr1sBhOpPzlws6LC1bnZss3OOfPU7A2gcpn7ioOMHFtO29lNRt8oIdHz51yjGTNYeYOshr
Pf+/4q8Qz4tYHxNy8xlT5+u8aytd4uwEC63bxTpYaiXaEl4WtioZF15JO6hkCxfyjnqyiF7s8x53
+Y6MDuGLixSPf3veBNN+tAWz81tUg1rArEQvdN3K7fYReTv+Hls0mD8Tws4SwADyesSS2CV9mtVX
WnvwsLn2QAtHXA5vcn2AI6Qil86S5Dj51MwoFgztic4fuzNmpXIPtKt2ur9FmScayNLULYGOgG0+
uh9ZiBg/pcdOjxjP+fXF1K/3lU3eLwO/2QJtncz0dtUaq1FWGAOdoDV3ePdvbdUHz68dRK2x8GG6
DCl3FZN1lqaWUiUjDDF1QmZstKyBIUDuIcfbxRJv6b/bnbry8USPFuYMwTKeokWHQtDBoKEQRCmV
07vz6tuqy2iF/8h30N7KHG8ak97OMPWkUPXr/T+mJYKlHMjCrWGIqUO/VFRIeY0xOQTshGnGW7kt
LrUqXoXJf7BM4RCtxgWxaBVlUQM4tx7hYUt+D3dg0I7/B/skEsq50PLSFAfsxWh222I89+z1weBT
bADYtcZUMKPzr3K6SMZNWKaAkrekCMlb6mqybBVsGgsmF7y1tWYZlVOrujMS++DI3x33vowuzzXu
wqaG6aHwZ/9p4Qv4CKkEqn59Jq0c6HI0AfWwzkV7VxRNHOeysta3NZKZApB5JbSNEtb/UuFRil1M
Qcd5hLgRlTlUrads+2aGhESHCfV8PSzZtrNcXwz8YEDJ5oqbSBCKzbIAXbcuOOJVwlzOk/rpY1cb
tzHQQUP4VF4g2OMgQ3gV1lN8dBgmL90vMuejVS4xFRXc+gLXhnxHvQohm1ufwhkY9li377oPZOxt
00HS9zxNey2MyMTH9p2jlX3h5A07pING0DrGjW70CM8KLLLx3Ky4LgZ2LQVi52gnL8PFQ+ywZxgr
S0S2tW72/Q/KdCHHCbRhZM124C6lHaphQ+JEPwKWXybwBkhd/kGOD8R3i1RiacYngzVkTrNFk59l
NUahXRgU+WAjA98KuBhWlQzY/5oz7lttEFCPn9Y3E53UKi+H/HgF4BHmO8V0QEEdbuBs/LFOTOvl
WsyMy/4cotjARW0hx30ZdYdEh5rmSuYbT+rcyYf3gb+AEnkuGmLqfUwI/aomdLs6pVnl/Z/+igRO
D3dJvB0TGzY86Ux/NSqTe5m6ftFwQ5Yx/C2prje4LivAzQXLsAM2yLMMXGi0MQ8nkG+1Gwqt49Uv
WbIy9PbULUxXThgKeFXlJ3w3ON0/OVjK/cmclraRnQJUw6/UrqN2KxI3pIGNOx22dzi/W3pUtnK/
CjFs5GLJ1Hm/DWsfdKbO0bXq2T6t+VAhGFzed8c+Yk0TRdr0EkmX1V1TsiGdZSZr/ci8xRvVz36M
7u7dM+1kUK41RBmV4jc1MCNXXpbYfkwdsLj1lEXekeHnVKk98pRfupi6S6ASqgxcCN+o/OyO9fkR
hWiv9tSWbNkShWfyRK5BqZf16EPSerZWp9z+v2UGtNUoKGwaaT6Ou0NbyPGVgYxFJFAHeBI7K0FK
mlB5/YoYL/3nYTaLBHxohtpldCFeaG4vUumsprHM28cwKP98Wpj4+Cf3W33Ew1jTEEB6FUzq3OVz
95EmJeR8LTIuSjl6Ux2kOGjhL4wVpIS4FG/3q44i36YYXYf+uVqMchZ22zAtA0v9BGwNAktuc8S5
4saIyhVO804yQVHjlfW/V3i7iRy7C+gdITuDYQtmoMxrcqGXKAIBmszn9ULWEmo0Nse93dZ5r3sK
UF3Gfa4dM5Y3zClZLJVDm6D2Ne0ubAYkLhD7W7bo2ogdJQNJKubjoSsXs8z3zrpMoEjD792OrP2M
/W7DyWFJa/6ccBqax3IjpXrWUOI3sT2FUQksdGF1aZF1P+Te/oiUBdN91eoUYOdanLnUX5a8kbvd
eFkVqYBlhzsl8pA3VVgq2B/We75f6upl92FT67+ztI8S8Ph+zIXzsgFKu5CQGWdJ4WE91Xk9lUuS
WSfhf7zLuDsj3OYI06kLDmKxefmawtYeBRv+/OjaeXI5kHccMlt+wHXUvfo9Lfhqnts9dyF8CnmA
Mu+3gj6FN73au89M9PE4IFuzBYQjBalR7Wb/1e+4aFGjcJ8vKMGn34Ls3ilwcCd9mOrj/lp4usVS
7rlHymjJaa3DHKZfNzbEMxkwJ+j6cOlmIvGrlhdVY29tPa1T6CCPwD4mhEQIO7yfNouEiElGHIO1
vV0Ct/PxYj360qnJnIV8+o8ehWyXghA+QO/2tdeRuvqf5/4dUdiqHhONbv8Q8ir3AZApvnJBRsAw
epjsHL6C1eV47EX+DMTBCNXYiPYqbGo0z/iG78c+mGUVfBKpO0AFktqki0lszKgQxCFdNlDSVU2F
ppmkMt6sngE/lDSAiV3rCX8RU1nRgxzSr2L8LnBNvLLZy1RTs3Aw1LqvkECUw5NAs3neDxbkb0Rn
/ZKUdRbctaVEcINQFOaonh7zJJYIakS67z4OTdT+wJNiWdjAPy+4kOoDnReLTDHLquJB7Q5pbRas
EBJrZaIGWj4cQuCZLpzfb9Hjm4ouxiUEJIVO6i3ufAR4JEC4G84q5Wzyj5O08Gj9P4xFxgT+slNm
ndAz6kogXsKFqLTfWpRChuzrH2PLKODnYjMYf6YGnZyqeEaQNxgWGWgvy1Ip8EIgqAh2YmJ4tHSe
kX/TmpgdlRw42ulF6LvIGRXUubjxfKr6d2rAgs0UngB8XWUSZg1xJ5GvVQHZGvlCBqrQbETuataJ
OUT1q2f+T/TQ0iQv87VJAZ7wPVvh0OEskFNtKHaqXpXkNoXPxS2Tq6N21YcoAYvz4NzBcoWDQPWx
kDQacbhwi9N+tLFse6fbQn85mmMRhUvN1+2x20QLbEhi0AfpqhiaBEu0rMhIVUijUwcMDhKCAzQd
yMkj0EquzYiPiyN5YcEeOiPjfLfowMpOZB71H6eEAaqsn0rXTAP44eCIZ23ZRzTtJYAmskCrQrob
XWVmp/0QtYkDmymK+a4siLML9WzOX5gCodOMKWchLCikckMbFwTc+eyBzfKAE7PQjsszkvVoXW2d
LA6D0fPsxcz8hOyXyfpMU+dWMtOeLyE23d3+pFThzAHrhsGwi8sxdZ3KfRCODy04pdyRXQyex/0N
BVFTFNS4WrSFzpB/pzwBxnl1m5hPb8xD2BhDYEyzK3x/2TV58sKxw7imthhg31yibBGi1PGs6M4R
o9XZXBCIJo+4VP0LA0adjj1TGdGkd9MARajPxNRaxlSmDOiH7javH+0YR26mYZeLbuwPjFhurRXz
cxwPPHqn6N65tsO0rpnwjtYcv2i2zsiZWTLnlp0Y9j6xaWUFUdjajaA+VfBjbQtWLeAqpQtF00Dz
D/MYPu3DFz00uWzrA2MQ9svizmQnUbmnP6t7VWzNdKKDVfU8eIOV+TqUP/U6v+9oerkRTyH6wrdf
8+H6VoyakuK5gXzzUkfaDh6iXoQDVD6GmDzx/QHUipsLwYLPL3dv27r/Kxa1bXUfK21rHeFNBOVK
/F67InsG2CS6olLckxF9D/Kh2On53FolMpItU8WL2ZVMAv68QRy1cBy03cP6gC9aGfs0MVkfg5g/
TX/z3qcnZEwWwwVtznE8J6cbrt2aXB2i+3GV5nHkLs+fulX5UyzopS2twvcQiPSpn3HvoeSIQbMg
h5Y9a3cTZlHN2X7npWF5DVAcs3Y2cAnKIhB52ADmnA7pUnCu/oE7Fus/VO8pqmzX/28eYW2bzSZp
0+Y3vXZOYnNjjuyEtffGJnwhqVcmZqmlskoctUhzq6gh6bWTofqUZkMINo1skFnCaryIIvUNJyxo
8nlsw1OVHnTTIMC5OSWjMoi3Np+8ApC/Jlcm4Ep3WaQVWzvk5CuahBoh6vt310swODKJCzGIA+T+
dWPpEo2fWq2fI4wONCoUP4cOIsGhbOEB+djVAs1zv7zpxUC9swZephDRYj3xtVelbFZ9mnVhpqfe
EdJ3nxpk2N2KuborEcUhhlSfiMkGd96rAnBPCAJXYzLR3BS/Xl2KDQpRODqhxNzL1jwXCQ7I4Q/S
wO+RvR8eUIBUEIL8212KaPk2yKDxK2nqUfc+kxt+A58IFycQZ0Zg4kkp0uch5XBSU0QR2dfSFV4f
OiNIjopbAgPmDrngFqyp1CamxAFrMYL10zeUD9koY1NNZfiWtnJ66emsBoV/SWkryh75ioTxRyuT
l2BM5zk6i1ilxopFkEl2OAWnDFkRwiOceMDI7cT5Qzi1EDfGUXQflFHGyyiF/kZmM/gIpYOJxdYc
Uc7twgGSeQzkiLnhYwZqZaqNKfUoeEBf8wwECBDEJmFxRzia73TjHiW6kyF8xUXLhFdX4ZXPYurs
yG7I96in66OJ0IDp+s77aEMZcC/kCJMm1uN1WM8BYPLvvnJ+4oAAqTwXjaaaE0oKIIFjbWkoi5Te
otStGQ6ePBsJICbhOeQPr5PZUV5itXj8tAGmIqpAiBoUL21GRE7kI/5DMEezLFVY0QVRYLcSDYqN
m66ImUcrfqZo62zBIZA4RL+RdwmDQLRuCc4sUgJL9nPub94TwYx1i8KLl35YlrlqI8JnxRg6ObQk
7L1Vjucfy3GWeGr9+I9io+6WiZ57EyeOYIj37mB5Y3AMOITiNvEmIoyEgVa62GblWDLN14KqEXiI
/y+oqDLQyMH3zZC/iaA8stMPR6uJeGU6hP2WoSSdgKIUa2sBGKBf1W3V/IMx6OY400BCFAHgB1pJ
MW6bz91k3aHONjFJlWOgek18hldSewUe6GGluf9xRI+5xZ0N/mUp6wiozdpFktZo+LIss9O/zmPt
LmcvIomm3ltf53zOu8K9NC1neHbcNTTw+G6z/ukM9lXIWeEDtnQvg8PkvID7aopWloa1pIz29+8V
zMimpj3VikvA22lJuCFQDLFOvjh3dtuhUeluV8LFuuZ1BjzwkTIFqfzE0QbiISVKeWpzUecLyzxw
8fRSD2GDBsYWMjKT6NlzZk4GODFD9tJE3sOFe4+jUqVCYNbmBRcRWRMny+qbtQeWUAkGS0/usri4
v9Tt1qw6FcdUqOhKygA82SfgPRxwuS784G9wZ2qcdU/I8P5wXxq7SCxyh2ngNLR+AFu2nNnLePan
MPwyKp9JNvBy3yVAJqEO4RLb0o53lN50Tv/uzvJy1cYXBD55UQqjTvsckabZ+uB1CUYrre27wtTm
2VYiIQQb/rVmhVZeshn/1NuGqnIMJQ+8npopodnWqIZ4AvQtIL552otkeMRw4oq3BfNDPggT1hAn
kCfOcO5yYb1GgI4xN7qVdHwiOjemOTRVdEf38UvOiJ2fry7Q0bXu+UbsbzA28jlJjtJsGtHnq+Wc
BkdZHQyew/1UnW1Ktcb1q6fwGzMHdGtYgDu5NRefdvQEqIQ71t/eYFY5NoIvdt5VNv+AV38DjW88
nzx8kcKaithNQO3uSvplt8lbpyFsGNkZ3NkwSz/ZHenisq2+hLZid3w2Mju9KyucJqVK8SDj3ELV
bhkhNPIL6ctXsdDKI/VRUcJVVVDSGQqchh8KDS0Tbz+UZMs9EEiMaLZxRTpeU5CctTdOuwhMDpHa
1B7rIF5/jukhG4RKNjSpn7ppy4wH88e8S79idCWUKJBLCFVpxqSmjKD1SKKEfdPpYHNC5gFF3k54
qkhrvqH9CCfNMWK6BpbTcE0pweOq4QdvDtQk3WVw5LEk6Vp1a++aWC4oQgtbceBBVG3dROj0RrpJ
zou8NPwvsE58cTD5Gw/gNPfcqmyZMqoShTJ6UQMznjNEO1tMkZ7t3H1rSZoL57ziVLvI7tPWazVm
R1vfmDoibVSCrbRrakanAnI5z3IT8HbzOI7ebJqV13goK9izoiD6n+JRQrH08zirj1BcFM/3AAZj
zIQKE41uft9oTEcWn5ndcXFdhfdHQj6zTIoT0st1aNM9sdZetI5RpSmOtcanzMVYLSWuxtduDmsS
PH91au56rMBjUgTSMcCYzObQxHUkCjSFKsAAcvs65vU1n18G2ART4W4Rmivh7C/iCIcZRlAr+brU
jqJEY8/KS1ZuNY8inCYTym01pcZKEjp+wpMsBWEDONgICmIfxW50Uxk0Kbk1EzX1Gi5vKIJ4Oojp
UOV0WVzvGt4oGIkvnHVzVCAJhuR8aqeE0DwC10qCWNXtreg/5SnxJ+AS9CTe19gbLDGTvc+FOGbc
APGN5yjWCRMW+CMy4R7zczD7nCY+A3PYU+qddLSZglWBMhOaLfz3qyo5HD+krXt4K/GzoIzZe9VT
5Iy6OcYJGMAl291vk3E/YlejoB81aKSnNa1zKGeenRXrL4j15lC7HJ2ti1q/mLhPoucwyyDXZEaR
VKmffqPIEbE9LOoJWgog72TcKDK15zRMS36RbFGq+jyweueEL9I+12kcxz0WH7Cq4PwsgXA3jH3W
0NvtIOM2FRPGKtasHgirE8YPXLiuoIg/z/A73vvg/VMbL8FuHfM10uuZb7B+0gtibBwIrmA/z70k
xyj8mYKZqlX9AKZfq8kS7Jn5g5kVQUYq+2hZ1OSnhS8XZQkFhPHiVx651mS5l+6a5mZ2We9rDLSq
c0rb6MFcBaIJs2FMDUMtsEEDIRHPM2dfpd8+3MFO8YER1eDmriXcAsq+825Zgrrfh8nHL/vLogt2
6TN5BAVwdQX0cgLnvo/07d/SMzUCOVcF/qm7LkWWOvY306Bop9+wUYjdHxMbQJQK0UfwFhzLP87I
VlPGUAFR8yqxU/TQEubSfn8w8hl7J/QQ55OVhzNgLetdklTFLFqVzxVRRhFa3VtGTDYiZPm1K7f8
FPIAM9+iFm3dRPfmwR4iQ46YHx9cuJ50sskgbyuzkYZK9vez0v2wgQ5WWxn5W4E6VdhEN0Wd1nQG
qBWZ4ZyVlIpzCcDqGrhzTCYYqshmV9yIUqvI6Ay8YnqWTSzsZaktbfiiFwkusjJ0idSQO8uuOmxm
dI6wFZn1ZgczEebMPic/duVuoi1ZunP/jBITsHLkR/eEXXrOZ7wTIfrccBVDSYAhkmEr8ixVMrBd
7ZvgY/zl0XORVp3RYSCtUICA0TejbwuV2JnWgdIQCdED9VXcVRpT7AMevy+eu9gCP6ihYacaL4/l
6wPIF5N87iC7RemILz8EFxIczMijR2qQ3OjHJmolVEwR5DA/O4uaFdHWX95mN0I8G+/8RQ0YHR8C
zsaECovJ7fhRQsisV8M3qftCsvY/4FB4zp42IYQx6oOUZzUZ5tE52Y4Z4FphO3l2P0/9c6OnDg9A
lFftMfbuYHRJ6kQVub/eTltIojVW98LJVX4g7qRbPA3rvuSla9ScOGpVYmC0AdsWVd4/LPdF0FJp
+jeiueRLhb1Gu+1bfeiqsNG4PjexLX9OLj9g4Fq7/AL8O4v9Sk5Z1IVTjR1I4f79KWS62RfKn/7z
GYHpi0uRfktrze2UHPvM6BzaIXmudCvE1iCOg8ysWdXNWAZhvBUxPEYxIPRRhiLUo+ZTsU5iHsnD
7gum1XihcdOHUFtajb8fe19L9BE1C42yof+0dPsyPXhyr1NXZpxMsdjP+KBG4c2SQI2UR6jg9x+G
9a7f78x5PJ4j7dJWUAsby3LHFfqaFPOIKqI1wUdl4LkkTpQ0sQ5jy/bktNysQI9pUQZLw/q9QpQU
jKePFRlUvS9lv1CJhD5hSaKrBl9SkxFRNIQdVdQ2xoXzHr7P8XGEDqC8kad39SXEVG2eYKGw2uxu
XB/1MCgF3fnjuuWBxZQUvbSz7o4VPa3CjFbWiXMC46zDEVnjBOpBcuOQl9r9+E8w+8s+DNua9Txe
KlAScsiPGd/VSk6YbVcXOuMGMUy+gVFupb7GuJOSoxKXPoG5k3rvFvF9zsue3ik0qlFH2f+xCmJc
mIdfUNrz0PqZ07DG9JQonFSNHVrjzEDinMDVBkarxfQ9GrS8Cqdxjj8XSg6VynYkeqiMJL4ubIY3
FK0rNqgoGirUZkIs21gRiRNjGgAZat3rLvhnDNglZSF/AGwsH4iA9BmAGoX9oBoJcprLaUni5PLY
IDMv4Elw8gZr+NnDx7Oh2PIgcAVkS1K3aGfNpMJdmAensnovN1399+Mi5rHvlGlWxnfBOPPGkA03
2J5iGeoBp/4BR2RF6zAtrls2B5MNPWfE2hFGdkFcF32sERDqrmp3RqjAcwNLELs/lFCgyM8sx0Ch
yZivKGufl+WetOMKjbzBw1kYy/fJWkcaJLjhLCe1mOTedTvmH7IYu7hQUwj9GNGVCXhOCtvzkXH2
jfrngpYz+wSpsgJof19Girptj+3zi6AlPiWuSwJMzjx3/1/UzE+8nJAZqBAKm2VPnQAO1uY9dTJN
7N4Ee6tDSPGDtTYMj/VE3e0yAkfPN/I6RgfBlHGykmzM/bTnKfZZY884TiCRYe2gc5DCTV9V1ajN
xQbwEJ+Unf2IfzQm0f+f79Ol/b0MN0EkQ50icqfDxWCAOtQndvi7IXUWgMVXaSZagnEEh6uK9CO9
aT5IItgcu/eSOPoeD0i9b3Az1kI8Q3EmoOW8Q1DQhldFaXBbZOie0dOctlnuXJZrI7N4j2DJ+WqY
sq7aETYJwp55dZLu+1CZFcN00ACFdARhuf1p61ulpolrZ2oJ6Cvwmz+Yegt6MfbDYj+nFrrk/b/h
xhimQ8G0hvnRhYnAmakjhbpgibSDHJg7Cceamo0N5lXGJSNKfuv/9yhzAEKzSIPTxQw+e5h7ZuG3
RR1Xh/uhGvrUSqDghzaxPixgtX02BiLPojnNfAty3l/uDvQXAJuug7ZKda5kKLtPNxsIMg1Fxq41
/uUigWi32sf7XrCBhx/gH1MY7gk+fROX1TX4qsj0vi+OAhkA0+eYbNafu81msueAGJZ8Y1+TcGXP
9+KuDm6CQG17GbVQvccE6JVA6ccv74xfLS7c04BiEIzL+A+Ft30lxfA0R75MDE2wB3im7senLWI3
zEya8FliBrZxTAcaT7Pj6XaPLGHZvfelDjkHOMIT5hEOzFxouxyLBBKbJ8dyCEVO0tKEIn85o8pI
5oO0nFnDE94cQhxfUo1xElAM5qDjai5jUbDn5hFJKx6Oi824QuQGElx/ZffVn61fKUO3fr6NemKj
0bwUFj2L33Oo2SiqfZsRKYvFobYyJRBQgz8CP2ZGLwZZerZzwmceXxOz/ST/33IHENAdK1tvE5rJ
Yl0KdwpmI3kBDJsthOaQkx+19lFbsxZ/r8RN5idIdgseQwPFTffcyNbCfAn6ioYpG8DgQTXvV0vP
jg1mm80bpgBZeGanl+mjzJ3xaGDiuIIjMhiTd620E2VBD0m52pvmKwfEyKrdYFINB4Z6EsXzMmfd
JPvkM+BwwgL2YhZQG0DNwkY1Cs1GLakezZc6HRL6A/wtpHkWUMQ7fFX/Gh2+yBd0jSbH+tFBsj2p
P3B4ej3OW4HHCzwk7rc6kjAisAoPkmDHfWiAV1cTAS/o0D3x++xGxkGv1seSiaxUYpUEXj6SG8O2
CwPS5bViHifBka2CqYYoot1G58uFTj6dLtSJcYpCeRwsc+wSAFzIMqvIW+V/GsLqU3VbhhUkXOGq
ee0/vWtjE9gA6wUTPyIyBWxy1HXopoXpsANemPEI5C/go0o+2Wg5IMR20x13miPRr6/jLzwMrLK3
Kvfh4kFIISHRd9d47Ye+MSUv+5HyAjBnEvtaHKWB6tIpP1bfuohG3LxXJxEt/5UwFJJ5CVM0E2+f
lMFshouKmRJt+K/uBo3Qu408M68E7o6C1FM0TEBRqVo9UtheaC9etnF1eLou2Vj2Q03J9FWRo+KZ
4x7vnUSahBA3ldMFOQowc1DFwvvwwKwuSneY+3ECWX88gbZJ8Wsmv7CdVuRKStyJQMSsv+fVhQai
9V0Eay4onhU/Lw1wL0Wpi/3xIXz3g036NlUJF2ny7jJTZxeYpfX3U37L4GClrfki0IqIeHUaKvxo
DjI7E4M2ztPKz5vkbZ67q++sNchTnVxq1gPr7MT/spFvZwnx6OQjz2UcKOGmc6WOqa1xeHkyRmxl
dziZHqhK/NH5M0nbO0E9/1Z+geONKHe27KLi5AQSb2pTEehKlKCcsX9MMmSI2swIroJXJhlKxmDK
7ohC1wxPbutpTu+9lzYVIA21YWa9/q3xPWSgtukwoku8GM6+D2sq/vLm2+JsbPdobkqxcMPuoSWo
BWK5nl5Xpkc3ubXCrMlJt2c9oiINcoXgAdyroGWCGGH1PqrAUfiG4r4mYxi73jXucXPg7F+16+Ns
nWvHWhPTEhtO+dtruc7xlBSXspG0Jpy7mp3GDRBXqx3M5U6bLIxiA8d772fGOU0C5Q1Vpa3uwUGh
sCKxAsInNam2e5gruUoY1uNYHHJJqpVjczTM1ECNvfc9F5kP5vt6uld1NVvUcdhTTRbhPkf40oaw
SYPlzNLGqZmx5xXpArBncJ4n7JfiXdfSabQlBmsWWjmtxnalSf7KcjjOLqCHlcNkiRV/GPv7Ltk/
J6AqgzNge4ZqhFL2pGGIYyk+ZJBNLHlM/Uqh5IwIEYZeIN3bDcOxSfgk/A7ST+utVH9NWzF/SARP
9VSqgtlN14LKv7wYv80H60Ywx3o4h/FY82s9WXe2YJxCCNPF3j0aFfqP59DdWrTF95AbvwwuSS4A
4PEEu0PS5q99SnCgfNe7TuSe2vtDEX7ThRSZLQ38ciNexkK5pJ1YS0JYky33inhlzye65tmnJrIN
vygEX+MdP6nxjdxK7oQhRTO2Ti+dQ5d8grSmOiDdvWwZEKXWAyNTokooFaaw1AUJ5H3B1bPAI52W
xrY6BYd+cHdl8VBihkQi8eJR3EtadenOvsXjaOmLMErDyWtOj1D5LE+C3qQVNRB8r7dQUWx0NnO1
DBixdT+vbVRHwJy9ldvMhKV3gzaMi9BTz/PfYZDF7udeb/jqLfiW34yNwpg22EyFUvFHzXtLVPUq
qoHBolUkSYZWpuhYyqqwLhQy40HA8d+HEZDshHgbY8UhQuiZY1SSxa+f45RUC5rnKk3JQWJmXhDS
5AyOwvrnyVincGZlBQdDvxzsQvK/KHMUt4/kOVPq2Kd5HpCahetF1BOuc1dLFe5j42Hf9rgLnwYY
Ou+LdJdXSZWzEBDI2oZEnN/sYzrXRB1BdaDqcOw4aydYQ+VaZr2TfLUmszscdHMvEb1YAeQSPzTH
kQS7uvIimy9PPLPZqAnfpXbHKco6p/ZDqOb2/OjV5ic+7YnPm+Ko9Usx0W4e6XgtzcHGELHoTm+T
rV77CSFdiyzqayBx3vM4BlQsS1XkR3ACJwRSMyEq6KB3hY/lhxdc/FLTZVcOT/FAB1DOY0C4tQ7K
YQUi7nmDOpnZFgLO2ukZd0PSebi5rkQ3Kp1yJ3jyVIA4+dW3pqYB5H8kH0OlbjHanFZlf8jDMsiz
mPGghKtSAWvA5KQCLTPZxxMnxnEn4PaKMypyCY2AzSqkcGul/5FII3oBa0QBskynQYk0pZJMkrll
X5xvoBm/DwtAhNCQOlqRXBrkmXSzEckVa35KhmnU3K3pouV1KTbPTEIeRtCQyF1mV4fRkLRidTr1
lgHch4IQSLBqfw+9b6KwvPku8EkSVAWsga+a/touFhN1ipCHZVukoRFc0zNLdkE6E7Ghx9T1KEiN
zGokQq8Dub7vzmdztiCEgKj1ZLAckR5pKom+QzJLjP14UvXULEevsSbL4JmJg3DfV0wkMGZ4TllJ
6/q92Vm0uDQK78Sg2+vlPvgs4wj7NmscjoRWc68WilJoboI0PPyKUSwcVrmJprhf0ur2Wo/+m9j3
GTKqAf/tBxpRwuFKhFESq1meH5wHy7KZjEn1xXmtwuevZag+xPduxNR41fez0PJP6Q23qEAiYEOA
s5e1Bd9NXyN8UkHe7emrKol0s+Kx3p0hKRGZbGqxnmPMSJkl19STMiuiVXMhTbuRv8Z858zivrOH
2AWQYkfEh0ioGh3qSq96NKYNcJGEhNawUjfnIdljZxl8rQCJ6OVg0Gv6gI3uBjbksua2WyU98MYp
3aXirR5gYP2qeLKQuZ7BgAT3f21ZDB7fcXU0NXxo6SmbDttIj2rv0ezPviyOwDxxp1bco1LXnu4r
aqZdXmXFT6Ns+LFfYQjtfghmBx1v8Cp/aIsScbsPt0IX9x8ImTZiMxyOFaMNqTggiVwNg8ZYvcbO
U1unwOqmxJFn1L4A7Cf7+vV2kghvPuABssQiEYxAZb3CIYT8OQCpU/Sb3siS7w9bDvwIh4Ohz/37
Uas3cCEXLU62ay+kC1aoxkzplg3dBl2zW/SzahUjAqTSN5m53NQMJhCrk9hDwBtXwSSDvQBFFQyD
W08HO3BdXR6iSuWkWq157f8uVk+gvkEs7YSrRpe7BernAxqC1cTztVsIdCex+QYKwqPCgrUxfLqz
4i8H+NMNIbk3/QlBxx9MSwdQJehZuFLQNHOb9vplb1pVtqZkgwnNcedwnof26+2cg8NmxPfoOc0u
pwCl+vE/NSNVFHWqVItlMHtOd2RrYXTUm+gAUgQr+6Cq/9rBGuYNJmBeElPwcpoGN7Z7iaFKtJ8f
Cx0aDkTjx/ASE9mXpuv1yXkq6Sxj1nvz4DnT3A8TOx9PNnhJH2Gex+ARdjHQLnd3vJlgOih+a2Rf
UMc+yfs9030UrEe5FDBxal72uBJSNJRbB0QXNY5ZdqYYqjjqMRg+zvkxdcEpFp41XhugdIscTlpv
zCuRaR2k5Qgv74Oo52uVJlSgAf6ltyHT9zuYq9Oud5ofyFf9+mb72rzPZZSV+rBrvTcKueRoEmN+
I6/+m0gGYrRrBsa6UVHAN2mEcXrxvvq7s4VsdC4ylfwIkXhFRVWl/XPXIBcsqNYwaPj+xwr4BA+Q
0irNA6J5Ffjq0/GtRXSlwdyG6ur+jV6eRw5qgr11IvlSpa7ZaJ66xGrB46T/TSsRl0on2qNA6lQD
LrT7RjhU3d4YUEodDG1EZeER0x9ioa1LFnixSNWMxbjbFzPg+/Hhkz7tptE8BmP7Ldmb/4xfmZeq
r7F/7GcDqHUiR1Wltl49XmhgTxgq0KwCqjEdkYInLHawMkqosUtpx/HE9JLGm2zjOdzpZGfAQJfP
jxiKP/69XtPB+v2RB6aoIBE30DOxh9NOYAr+P2Z2ffToUCMJxGx5/gd9HO6t0yUMiOSSL5ERL9vP
jDHqZS2ySkzT6+LyuYoVQ0ObP8UxL+L+5ucpOBxGfRkpOyJHPsH3KqgWxvDp/VOKrqoqGDVAJu2O
AXy4NePnAI3Qukh3L3J8zanw8A3nbBZF6N2FSvCEj+tMxzEZq+XZ2q7J5svOAdEQ5E+pd8NtQMmB
yqslPLFp6RT39F2/JN2Tx0EQtvItSZY+cFAB4LayhOvBoQFxYzYvt5N4rhJrVxwWj5nbGKV05/iH
fNzDcyn1IhrHUQHLHyF6oqEZrCoCT0seGhu0ZwwRu83OO92CLCVzs8lGmn37gJdmBNasOG8nIJky
VfGkSc7ZDyLmO9O2SE/TNmMGc5vxRASddIzFlwyXS51ZwRq5+6NqKE8ovzVxyc1UjNN0ni676Ftr
hZJLxZSOHFQnujnu5wdBD+BjlEUnSdbK6+/6q1YWlJoHCQ+DMYKZlkrtTV6yzTBFenigvu/dO3EB
OZH9dHOrtNg6kb+zjUxwA6x/SvIykLpCO1bQPYNX6UfLZZSSPuRVcHHDbi0f5J0kSUcFKEVQJpGs
xiFR8FYguHMrcKIqAbFCwXtmllf6821iFe1Bidr56d7qpxnGhyOwueO0Rm/461RDEB2mc8uPDk2f
8hYsQ2at2HAMm0TVw7mOk+JUXTYa8IZS3o2dRwhNWeCaaM/kETsjStSwuqidXTYmM15w9J+O2pjY
B/08WSNAJ9Qyr7w6vwG9KjhWcSRVXEUbqjncz3T+e+I3FS9lvIf3AeVx+BcR/nq8y29sc9eLO8Oz
lv87UiMO6t7vX/6acqsyCU6Ets3KArzGspEEd9IFmPrO4stWh8sNwouqLdhwTvBjazNCCqtID1iv
eLgqJfWboNsDuutEuX7S7ZYxT0mubCY+d/qpKVEQQGJyHn5dF+W1HPRVy23wl7bWt44Oc10oKgj5
XqOWf9pvZyOVN93F8Ww0qHDRlYnUunRT15O3iJMszPgtKTUlAq853H2meDayvPDiDkJuRG5Y91e1
RQZzn5JJUzUvcsOxAuv+xfajIs1HcRpW8bODyu7vpuxSW5CpXe3EcdDUaZw0nbwt78OT7Ov22hrZ
l67cErAP9fz1CBI2eHxR5WClhXDH0c0Cf3jHpDfjlbUYhKBYivpGG1juFAv70PJ2UkdbMWkkpDTx
wR49Qo7AOpJ/QbjOSs8NaQLXiD3IdZ/iiOchCD++Zt4TiFCPYQWDpeGfcYitNeYOBLR+QlDwQ3lC
AAF7FpEcYPG9AVx+qn5joXCNk6t4x7LLk/pxmyZC5hwuRxhmwAMohWjSJOJ21vlVZSufv3V2zAPq
f6hDLlZQvL6PGWi3wsjqozIgMzOp29l/P1cxgk+AZEeFSGwQ96MuXA5or6Ly0IEj8Pj5pMuk1poz
2NWHaUqLPMpnwp1mJ+B+WVeOShkaNQqVw7i6nbQ1bY1uHbVfk9/z4+x152SQoDxLiDToirLXlG3V
ZQSVLfUmwVBuPOQQDoaI0ydTyvGsJAvQ88X/hFIaaqr+760t/vqNX/LbhQ6g52lT9s3mIezClZmx
NZCO1BkCu3swvmKuXqZKum7nsD2A27ABnNIvRQCyKy+vSjAxpTbXbcYyj+ap4TsW/de4lFVqsCmD
Nvx5pfyxUV4Lgx0CGbQSMpQputxvXXqtNKv64PO0akduIdjGjXsKqQdVi8KP7laKRaPW4uVEapD3
gby2Fd+9LJRhI1ex4bidMSFuqB44GPqfAoe6vQsLjHytTcHjDvimB9t499bGoma4049ozLC3YNKr
8OCiAPDdauuz8NlNTeg2+f68BcBdLltCGBC49kWuJr+2jW36Nw0D/59jmZUPLhWImSrm5jQRzXcu
t5hkmOVUnly8sKVa3eO2JlTNnvCV8uMkMKE7qTPHV9dNXvCrzW5+DBqy2kXr/kQPiCrAvazn3itQ
7vu56hkY8FR926ZTjoHBwpDPvBVDXLSBCsimKIYmtrYHW7acjAJOPGp8+n+6VAk69UYyKW16jWBx
HTKh5wZ2mkm8WYq+nmVi8mP57Lm93CNqQPapKqPyHgsBQu5fqQhgqB8oWeewd7k0ler1ywlYyBiy
uHV2Da53keJ5MMN0OouXsvBkv94Pq6nDmXeynQdRiduNYDfh7hm6nHUx2uBbzcxztZOk/bC+DEpJ
4wCmLkaeRvT6sLeE/2tBJUPppRCcruZZQkLTsu09hpT5Elvd2zSL6r0+xY5gUqiykPsQ3A2NDFz5
rLEEygsBymV56SJ6TyVkGiRZnbuWwlMDZnc/w6xMH20HDDwp1VoaTkJcBRDIzUmtAaH0bt4KZd1d
n99fatoypA9TZAyvKlfEYYj6JkkzBOVoybAIP+NXrNwZmCMhttOKSH0RI5bEp2pg0rXmKqJOnrir
ovWceZtZtFx34uyTV5zT5Wn156HjXS6bxEm/0TQf2Ql/Th4D3IXTiNqOMJ/m+/bm7TyWxKzzRo/s
JLpU81f2eqnkHH3Wle9y9ZQYScfyU6Hzopy7gyjLTS2ElxH9HSRuJGwEK0u7DWdVsw31v46RSn3g
FDOTuVDb/94TUFdDZUQQ7srfOtbg7K85UuQolgkQq0TJaWqVz2gPdfackSAsIMya+2ufeTq/yVAd
ou0+r4/ULG9hUVYcMPdZ5dp9sxI3UctfRdyzMF0ugvlpupD7uFCsMOCZhGP8hAA7Bo3DaHLfZSrw
jereoKSC9T9RRdHyWwUZFlxV+ZX3CwcKpyozButb/4FTPkyrs0I3hzINH225INklafaZWG1SdI9h
onoRRZVe+iC8eWiRLdcs8y9NZwwKJKWIriZTRsTCsRF6I2FCW7Xf75xK1WRsj+7UrsQjNE5O+Mam
StsRKcAsbtKRf5L5H3MeSOy187HZujVVtNdh5XE+79qUyfs/9EVTuGz/PGAuaJaa22j5RoQ6fuws
2OHHWfqK+tsp+ogCuSmQeuD1b6T8wNXN7x0mY3JZiwPFhlynYKrCZUEt1CpG2K3TgFofisURXGR3
ZCExVlNI97bL+w57ldaR6uiNs48zk510IDLZupPfCxboAyOuZL2HjuwPnWO9QbD1fxacX+VX9J2Y
L9PrlHO13Klmzf4YbdNufEr8ZfLwJCOU8Pcx3COO6mHXPel5eEtnXSuB/jOsLUq6qMz5r3a+I4Ik
syFBBqIMY8mDGaE3kW3cOzy3G5zoHE6Yspy7UGGbt2w4bz+qil5PpodbC2ooviWDqxjKbYpqL8Gn
1QR/Te1ffyERI5Yb1Vjlg9/9cxu5fo6D5dnR3Stf0VIXGgFk1YOw+7ka8DHuW3WXgx2WiKG5QWY5
+LlcQTPY8jGBJJ+4Zl1858blmwjKdpaATzQv6nYGCXALYheTIXqsF2fDgHah1zlpusSes7yb8Tqm
jMq+Nn2Tu+pMPexFHas/Bpi4mBCuz7nvaiamwvtzuSIEwVXNHU+1aJf2EkRvNsL89QO7d8bWQ2xV
SoKTO3Ixm2EfHcy+/1GeZkkE2jFPq8zWVtW/5hkCupc8FKSLAR01vtDftpn0gldg2s+tocDzIT5I
vpiwVBiK90t/b29XB/pKRdioy/TCgujqgcDueJYhI+VyGhuOlQV7oIrDpg8fpNErUfy1JPu0ID3d
tINy7vIeD3hthprOkI4hOR9VJb8Xl+/VpPBC98i84WFMdMu3inTYcvX/QqftXOBiy5BdY0SHx1Ek
APIHTy071CbGWblLLHjbVbfKafydzaN88d1N5z5HiAIPVDgNX42Bbts/KRLaQmNzA7qzFl70ZClo
fvM3FVGHaCfWozn+pPqb0CRkNiHTHbkSsjlRiMu33xNeOoT7n+js/aXJI461PcK8ktrsSw/88nAU
ycYkA9X9s/Xt1wKpF2Kgq+PUI+OmLJV/tdCELObVKsJXo/M9Izt2Yw24Y4EFSsN1qJmvZhesSSFT
VdQYFlmMeFwjnJCO0AY3Xors1PYh1I1LzKrodWkfw0n4PaTDd2ANeRZOtTM9uPHjDHUigOMlxB8J
VrE1kYdktutCf9JtXcaEHsIiTSj66bOjaozbm/Gy1ZURAK2mFP/Ri58m8YI9ZUE/LH6aLNSAaWDZ
VRtNobINgjW0GI13qA2zZoCcgd6eMd8xDNeMnQeO0m/iqJ+mZfrBqcrOYzCX7VEuCi2vjpRN/ski
WnYqkRrTItdQdYll4Mm+Ew1tZEnO+Zwnj/B/+oivGAlxLmmHYXRHSw8D7CMoDKGlETRpmZQZOSsW
7fSuMuOVoIFl0fy2vlTQsiIiEJ+tbNUsMkHptUK9jykCZsbwf5nU0Xe7kyf/hkXYOI1xktiClzCK
Mi3JO741J1Xe44nOXmdH+JBjiFMjVtMrV2ZZRez0+Ib6YyLwgKL0FKMF7tz3C3U0RUgA+5/xEpgR
MH64HczVB8feBXJA2arn4HKuhXnf/9H/ahiqN5kHoIl93Qmh6jToDBo5QsdeRZKeLyAuFS7hKbWg
LE33VeSyh8kAtjOoKcvKD7by38o5m7s0Ludfcs+JRX9cyLyHJwQRoQMzhRiQoQDBxkCEbmnZKV/h
9oc/yAuswbRxaQ949nEGslQolqRKqftslFHTK5Eo4DIFGmV7GAuKb1Nwxrdi33pCGTu2ov8Fm7S8
gWm5ddhsiDq5opFxoeDsmFDWXfK6Ol2F1QGRV7JpHfDkRNvOg8BfZ9gNHW+tsKznLrJb1Tqt5iza
8sZ3FiEnEuYr7K7XyK3RC8rExsUojfsY/wxpY1i/W9+XUaiMkUjbzc8G6/dgsLPeEBOfG6Negvf4
zZfSjxT7BjWrVoyXYm6ZphTbsrAwUnrn9461t9+Ur7220/pMwzdlfx8XxJhSKMV391pfxCVXFXdY
1dJCHiBx5KrcaKS7wd+l4M/YNZksHNuhVWiUe25gq6OBHKK9ZyWR7BsvXFVhU5i3U97ZWH166lgP
sEE1T8d5efwGdtlNETksBcqejIuRD3kt1vNUM/HjyhUoEbp3JjITK7qrEsDkkl9FtBKm4plGyd/o
Up54FnVysKadeqOpALg1JbSXUjWz7nvdslneU0GAzogn64TJK4ibGVcphlKutN68suQQAgPrYuaP
ZT8e5T0gY7o3HSIEMJ0bOkXqrxN/XgBmtzZq+P3sRfaPDl6c1zHRVjMQANJ92W5lPX7eG4e1IbwH
QUqGiKl9k3EQw+uWbv1k1yx0jujY5Mf34Y5XH0FVDU6F+kt5zorDgBnukZYbrrJUWghEakNPgYok
14yu1YFEtRgSBgM9xw1hX29TXd0ekKKTXJHE8gXPcAOVdlyIDYcF3Pdyq3oDQJdC5n+EF+aU55hP
M9Bhr7ZQvMh/Hr1p4JpzeIj49ODOcuC2vuKIHD3uVtsNnQwRpdd/D4qYhvq26Sxe2xfd4d5eHseN
3aIaufwtIc6z36FlWcaVrDkmN9/bIf2HNJZiSkVk2cDDlJ8JLS6jXaA/D1ZvG26ePBdSy4OHlo48
hm/4qj2zx9fl4Qutfic+UumUbW6kzf7ebFISzVU1qO3F+8XOAldFNE+BvCJHJDaXx2PShZZZCfCO
pQiTp5xS0KPA8tGAdQdAEJvlaZXxbxfs3ws4+vYIimkK9k352iDcPGEsU4lXxFrRvnXyXgno+6x+
1k2qIeXLcY1xulbZTRMSjU+IcGxGBeJawlWGKvIoKg7IWISZFo/BQOu7UWGhiHSgF9RMSPdK5YBF
AKCU7UR/Zh+s96u5H4ObnjlOntLQ/qVcAQDMZxvAFZq5CyaGTxfY1MjnJmjxuLJK/G0fZx+ulBJe
JLNmj0FloS+4BWjzuALAEcB18O0QSYEeDEK/Pgvi4MMGOpaXU9Q3Af6yvtkEQVFFCg036/XmGTN0
sQO2eci9zFR9NoIqS8bzNJzLAs7sv47VEjLVXOaTKqj86xRW7M39ORFGImZBLdOUGMXru70PEaBv
Ja65KOSZP+4M4A4yQF0nDekE+rWw7R4r6hT9eQTgcB4wnuQfGiXZWI6HSnMmeL4MK+L7hV6wAgyP
pfsyiuzYEZ6srtPUQPrmL0hBPgUE6msj8W4Edw5c+mqByXTyyCMKfisJcyuG8vPWy+fVSDtp5JqC
UWwsK5u/t7mgCg3CQUw7c0ZTeJt6qja8DZrIj8cXKERpa7Zy2k/IaICO9lOO52dWZsrlJqoaKmHX
A8LzQ/cZtYNgcfjJn28cTfXeu1yv6RK+IyctkPFugsRKiAezyyFciYUAI+o7bIwwIts0leTNNXU5
iaMK0jYEt00vvfcG9KNy5goUcgfn1hEJDu6kDYzANVQXPff6khTimpOdWvGfexbUD+CLSqqR+VzV
gfbHbSLJQtutu2qYxPb2gcdi0e3Riu6fnNZ6hC7EZVmtC3chdFeUicVQFHsMVVbo43V/IcTiYnUI
RSMh4edlo4mGM97Qu/8gjh8OFEYEf3mwIhXnqmApxqDhYCyVfnqpTUa6YnrDmGXUcBATSZ1+kQs3
VwpFIvjiyTpem+R6HXSTYo9weYeyzcQOJsy3jJ1z9uhy7Abw128ZiA1Lj8c4TqeISybds2pl12Wm
/vDAFvFF+kwsVqkpd7aE5aktgsMjBvavRuKWvTU31AOpEUP4Sh6qifQnxhHEasLIIwHHBDervgPk
E6vUHrIm5MMMIH2T0Q/h27G6PG1qBgAvIk1lJcVw1CjqqHaBzvZ7b5MhBdFuPwN3krl0vR1LSJsd
dKc3waWnXvW5uHsmhiwLatNbK8aKu/qvkU1OHfOszt31jBYX+/0bm4pg4JbWzzWaRiKlYn46DR5a
f9gPuKsBIYJ44v6op9rjkwHDWb0kQfe/gUp8mfkupdNzvHX7+7fkSZ9csOdmBsokP2Gp48YvRdND
tvwoRT21XhwiE/Bu2ebxKAGIjM95z6fs1WLmiEDHEvFPn5MOMi7qT0s01j+dBAzKiS4j3X6qtGpP
6kzX5Kpuc4aptZPtus6IzJxXG7fiI0HADRh2SAm1TN9UJpcicW7tUus9JwJGYE8wMoP+zcDF5x23
JJXYugwdnnAhvRzd4jgcegL8X6+BlSDMuUthuda1fHk5pgqFq/J1oKGWs6+xgfQpjnUF3LsBAfxG
E/UbZWwBYdymnn2i9YSifsh50mkrRfIlGlTK+mhHwUzId9NHsyvIt4PP5wI3NIeg/palAwhqXPU9
GDiugRdpVIwA1ZBD3j2fZnesupI/PJJwOiU8Ndzj4kaQCGvgq5lnD3Oec/xXkHCyRzWuy79yYjqx
W1Ah/Da8kDJs1SxroB90UxfXswJS6q+P1Ls7Z9lFkaUF3REOYDxlGHSTU5aQXg+IR6/GBo/KiL/K
wt/G//Bp47ZGwqHRJ0m11lhnCJortnjJkSJShvhHD5ltnC1Ar62mIraNgSYZvc20W2E9CZHezuG2
OnY8BgVkYM45mNHmq3AUV3X5L2uQB7Bf1MNogmcqL74e9z6HEBeuJ9PSCaCB8QJA7mx/E64AgFay
nBKqE4vCtwdk0NAWfNQg4PTqEVBxaMfEG9Nze7+c1b3cOkec157vpxVPAU1qDQgiZD0BlqzLwx2p
Ma3usqEhImz7JunDE57PaMzF+ZPSUOCqxCsjwHoEyiVptLswX988Itte14hxRhmPh3bmq/Ex9zBT
DTTSVI3v81dSZXZZn+QGgIlDHWRSigX19IcTk39CUy2MQPRpaNbaGSGerfpSzgbYcn2/EZ4sm+P2
taSSB43MwwQXDzsbFlSSxHufOL2VbrzbckYsDYq2m3SkkcgA6DPRFPoLVFV9NLhLpv4UDn5pkRuD
rxCzQHL1noa/tHpQitYGh/kaOErFFOmP6euhuMN5H7rYCOXX+EQHsTXYfWcN1pZz9a+yqAHryiQB
o9SxReQiVj3dIRfUpeu7PGbD16H5XB5cZq7aekI/f+IRqxoagmZ+WZJ9262z3zXca24vCqvN+VhO
+1WAVUy84vfq9lJzhOOH4DKjBsAo39qrBCYlrGPkdZi8TQo7ncAL1NRVOeLNzT6LJOLVdAqnpQIA
7v7jrVkcqnHibwTvCkM6SBWTsQXHHW1hAX/18OwC/paxcgszlcX3KmW1BPbz8v1SZCebEMjDdxz9
UpfckoQfoMxLLGMi3RGWz26bsFad3FvybuM+g3xfmWLUmWUU2YcIoKw4pMpLx45nkAZOXKOv/76R
4bSSeEwTYRKFvkfvFBLnkPyJQNFP9aXSlCPAwJzddm626vwjK7AnN7J7vLyeizI21yIjmLHLojNf
KG3ORH+Ap+afQur4KeLi7jXz0XUGR9LydRu51Wgc3RzwgIXzrAUmkMGI/EFuWbleuMRe9HmZDGEH
rcjghCp9KeNm8I+evWceHYWCLSr9mYslb8/SuEXue0EbiWgUL2gxtmAYX3EicP2gA5yKHvTvIQMq
dEKZuTBqw1nTSdq/ZBX6981h8DsIG8jt6xFW9MjiieZDWpVy8MiQjV4TuEyv20/WFlip2qswfScL
Ika9i7BnGjx/fsHJHdnq8ru6WZ+4eJttXy4qWdN9q3rMtkHwcpZ9fX1bt6KfFpLwlIHFL/Xjg/Je
RLBM5lMKDKaUniaXILqcoRKsvC/dJ9ZOAV/plETZjJx4EjnGEChy4ozJdvpceYYfUeaQTTxDRFV1
YjDNtqdSjXRVi4nN9VskuFKLo7m9ejfj0F2odglG7/Gw22KDGpagsIzoe1ANjJvDD1uMxno/XQgA
DKfMJl1OWsQs8KBJtCISGibeawcUhBCtxZJNvdfS+OAB1b/PNLFWwDdN4b142sB1oYAQrq7skNEC
HNHyoBeooV8pjcfpCZl4bQSrTSMJYDlCsRmlsVTS/RasqkD+2MwlNqe9h06voZcnowaHo/zMUfy+
CvMIV5/kdWwZ6jRgMOQ0dmi3Mwdbh6xWMYPzVgWcJGLX5s1ZeZ3VDgafs0Dct0Dh5LbvItTAb3/K
5WVe7pQkRKRF3EtKwRJngXbtMugYr/AsmYRwt/dqGGs7pn/645vxXvKxUmCYHrTrxogRLXMlMt97
IqORLe+nDu3oNGcQBv7Xzl5hxj13OnOQfqybVO4jvl3fL7wn2nqfReFEH2m50in3So9fIX1hVq6h
hBgEEz/aQ2uwbx5bDXMSL2A01fhO/4LQhnipgSrk8MCMkY4XUMhm0D7zEKsxEL2UDOpZjVVfv1nh
vhY7+Phfug/Ux6S902yQEdLBhQc5Vr/pfWU6Ui+LSlN6aifRIG5mhRirZeWcjUmwoEiZyHQ9IPuz
zRbhvajSGguIFgi4razYBHtU4z1Z7rXYL+MdO8hUKhTVeIBl6KnBXuOlm49ys8YhUTbXAuH4F2AB
t2mlwe+6bNvZp51aKUmC+LGEYuwB5ulJVeyUtvfUHCpZzn2w9vvovDCv0YtZAxeFak2bpvQ2YCRJ
MM20LpJ/B2xeNQF/5soaFJ2BW1ssjfFURmmmFfEeblEI/c7BOyWvQI2OBAgJeEKpBQIYm1V5bKf2
zFioKWFqp2co+gtkTeXRmCKEpZzOjUO/AKIcGHngAm4jXiLFYaVTBuZmRzSjmqQLNbsXy6Jh/oME
Xzb3Sc4iM2Wx8W1+qwXv+Wu6LjV2WvuHlBZp3uoCbqDAE9WdkfTpSHsChH8RAPA4KczQWC8xhaNL
7Xou5rCfGb8kPAzi4XtlM22c/pjsIwsfnptz1Q0+Wda5WCpp4yXJUf828VLbpzgXJzp6Wk6mBoO/
dSUIYTn2P7Sa/5J/Xajpj1yA+zZ1so/gcw4z0t97hkG3D+XAWQpymIWRACzmg+KPQBo3x9htJP3V
oaIDzNTN0Tvug/zFdKEl9ud8ywY5V1nAXNE73bZAjSAtovlCNNk24Jl1RTuofqa+p0HbH21y62Ak
6H8DQdVVF8WLhjHVvwbn+ctn0LPOjYISJQGP80IxZQg9cRU55c6f5eTFzBeT/LZIefeXUcqD+7si
va9NoBteLL99feOfj3SPayLLYMhVtR5DSyEVDzFLRV9uPYbA1W6vdFj08Xp2eA0MBPodLbA9JIdn
I0OT6iZdvNNuWKZxxawHqmohVSz7y+4OpLoPBfCz/QJB8cB3zuz2DCnLCO6O62evGVtkQLBmf/Hc
hG1wgMnJEKUDumAdEF5SO1fRWefuPlG2VhVwRAJBsZAwRkq2F8DTMNbFrfiTOw+RCRTCv72XCQP4
7uN9MbyHrZG5xrqPz6oSMV4QXkUlfuuPOjWOGOIaaBqvXtqVeXRhiwBvFQ0fvO6698WX+19h0TE2
Y0r75BEof0srGqM3UWz4yCDFI3kAZ1mAyNM9mDYIfaTti85VU10BIwAeJis0PvWpUyE/sV8sTYfB
H5yr2R2k5eAe+MDZGUjkCWu4q6uY4xynOUv+Mrc4Dsm5IbCsYvutDDl8c0nWMYcIgr+rCmH9R4UL
ijxD2L3Ik1g0EI4Z4TeZcHKMJMyWXAZ7CGc2B93azqitaSwzb0qlu9ONE/NGN8hPp3n0y5WnwMgq
mdSwmswgUYwiRqlwfIOyjrlH/o1ycmH6Nzj2plBy2OikOpU2RkrDd9Qv7b6CxQ4NlSXcx2dLxz+/
Pg7/OAYGvxe3yf1IngXCKOLR9QiqIQ1GTOEFWbpHOqzVMReOvPxslbJYrubi21hOCBQ2jdX55SgR
3OmPQvdkLRb5gFUvbCOmosp1Hy6OJO7drpccBpNY+N+o0tRJRfA3cPG7UKW/Q1HERp05Ib3gbhRk
ZJdWWHDGKbfMs5r77L8XSLAhySf9mqzEXR87dMziRmv+6AQzv5gSX0+3q6EtHNZ9NC7AL72xtS0m
eTzisGiZ6viYDOT5DZChl5YCq7HvFjtorLCTGB9OZjMUn0Nn2IxLksdCUYZZK0zzS6wJoTIe6Us6
ZlZ0tEYjC9U5OQiWHb0u5ojKE2j07fgVWrVMOCbknHsIyDL3LjCvS4JUubyC66tRPYEzpf68YNqw
AVH8byqHZDyL+/zn3r5i77A+1hyOCdK/uPKbOOXAvTagQ2kX4EKTDsrgs6lUE5FXhIh+4MoVo6jL
u5Px6L+8ptyOf1TqhCAQsuqHLhXwAKiQcf01AJZGWQ7u3Pwz5Ch8KjC98T+CWhIh8We7aALNbey0
VEtPkLbHnsp3xuuHgl4OCLtKfc7+aqtkMvI5kyKcCxeOzQ6urtDUVGyHh1mUl5pSPBL7TkBxv5l2
+UlLZU/nCBhLvZCk3412YHLpNQ/gch6kFB1FZ/2iuklOIboofCzac0T6MWzG7saadmdqyX9QY/wr
alc5FoX9lfjBtdGoI/ypG+cTyuJHnrTbHN8k/vMoQ0KfBrUvQo713QkoxU+m9HUvVGdG2zUrH3yo
IA1PK9DIh/0Azr/HeNapyap+Xwd2ULzTgMsGJ9H8hU+yZ9Ml02wi8LMSGBocGVr9fTGZAsrFCUtd
+XkXH87bmP3RQ8tyZB23pASU6qXvG/FAzPkHVtkcaB0HSzxgEvcaqNZc9XCPLsMY5K3iLeGtb0gc
8n9NXuj8jYvCFudDcCcXcL8BCSlf6VGe3HLPj4X9vr+sL3FUR9Bez5BrMZFZR1zukZMdFy5eKMtV
baathKHE+qGC9bTL/70zc4F/LMVHzLqunamtq2L91XD6BJ/JlDFqLGFMruOBH5by06tAZUCBRWaB
oE9sOO1EfeWaXPc3KFufqg0Yksj+Vq5ONqbuqFnDneI92g02npIwUwTr1N35vOMohiHZvsT2HJF0
wrpZ8/COglgzixrNNTis+gGXluIboJ/gBwf5zOgOVSCELuaFN/8zv1VwEl51hi76re6ow6lT4BJl
n63FxGepyOHjLHb0mZ1ewdfLFYiqdacRhaoakljpgaKFoou9jCKKJEtvLC2wQ9WE5cuUN2DOJdy6
z0LZctc9ELMfU3t6eTopPHY7ltK01ZZRfELcRbjeAi9KYeFQFYgWEDPPBsH0lkFqce3Mj+K9trli
Ko5GAK6RslZ1q4ZNVLztW2/YAnvq40iPBx9aAHaOHjgX1YTZZu3C+us8M/8zUGKfZuM1IaksV9Q7
ZBkErwgMZ1HwfIUSfeQl8Y0vWbggFG0rRvo9nDDivXQFt7DgDyhWbKWrkzSoRSgtZbDXPU6twikM
ig0cd5ye0VhmPuTRnYKZKPsu3AUcfma5We4nWqYoOLpqYPIitln5NyeOqScv96EWMi3w+ujK7Mwd
LB106+eSLotoTDzHSx6mewovQ4Cp03/cYhHPjBxEeoqPkAs7JQ9CixqKX1GOm6tbagxRbDy4tFiu
BmbJQ1N3/9dIodsJblRvlRhbK0VBvRc0OaSeh0YBOUMOs1iCq3y5ZTD7MnZi1FT7ZsEp5iBWM2pd
NJs3eY56Irv2JiPDYgjGA88zUTTlqmLeDEGINl7RlvV0oKm17rCREf3a4UcSI4Miyn75kKiub/QP
M5Nf6STetkIoWGJp8aGl5msrP7Nv5oND7T8FL4ykqkWU4GS7gkYrTfW33tLzQ6/wWAWThTqON0Ur
pdhw82QvawkiSyRrToj7hgNvJ9aGZ0+vv5WG83Qg3DcGKAI0m7sTSPINf9cnNcmBtu2XbgBVMlve
yWNDefo5hmiEu2zq19FHv/Md9OjlRC87h83Ma95XnfxIIvZgVK4xZaVJCs2kPrnJSxrySBYI1keW
iRMZ+STAgtpAd5VucWNar0Es7Kvc2XEF07ps82j6yWBye/unMa7Hhbz0O4aFMGBbF3iFDLcQCU+G
Eul1hQYimYFRbastQwz0na4kuMgSSU13O1FEmgl0IUrAOZOZ+uV06KWzmHnC3Y7EaxlJO3sY4ZWC
08jwOU/3jRJxsM5RpuqIQ8DJPjfODQjK7AsT9HwyymDm8IbBwla2E31ElmhsPFfG9CnIWGrNB+Q4
7Bp5JWaNrOgsECNlJ3PdmeQDtPIvNOkzulvEUD2BN4/u4TEt8785FMKCE5ddI1C0NXzGVeFy177A
BhcZHHUMkh8n3w4SDvigzN+TCFuKht4rCmBrSyX1urLlFXThSjj0AmYrRdre+dfaRbf5oEH48hmf
QTZpL6k9cS1RLM10eYw9fJ5YrZRLXhaw7IhVSacsQhnv1GCLDtTlxmPJDNT41JEVie6uCfffqW9M
QDGARivVnHaeZOAbID9o1BDX1c8bSiOVtOTCF74BgLzvIqEwPrecH8MoNZkZJ2PXgtIo+STiv/ad
TsXhM2WekO55Rhqkj4CXTohLTX7y967bcEV/GCXZAcSkDIgLdw/chcifxT36TA4T1Lhwq6axyLm7
ZpLwDru0FQ09R8szO9Fo7+Kb1INNH0TBfTHmW2YD7E0UXKoJAU+SV6D0rD42I2wx0wfk91Evy0gl
l3hDCGJkd25bh5k2GKyp18qjvgRVlP8tx6LZLUYfr8uF7SLZ1SIE8LGOyWSUTPCCKiycT5I976lo
dtguX3tQ50vAQfQYomz5A0gOZUV+5NZPoE5UF5+7jZVLIg9INQTaLN7bnLAv/owMh8oqiWkv3Y0f
qx+PB702GNiKrfBAgwqznDh4Gury0vZgiILBSJUfWHqGOnQzf0SM+AGDae19l0vhoEzuXY2CpfVJ
d3qgz95+iv3fG6Sv38ejA7Knz2riktwTxb1tTCg5NyoFDj324qRwyd0WETFNF+91qQZba1bLyMwM
NV0iEk4r2jlzMgJ42KrXhCetlbqLRsNJ/G/SEfIV1XtQ2ZxO6yXETBbu4uL633Q3Ck72X/UwDeSz
yk135B+/bW+sGeP8mTm45QnUxErXCcq1/1rWW7yoBlmXszAnQjhINDR3dGyff5BQwyEa28AoJcvv
Ko27XrbDxf6g66c9aczkZxY3YgJ3WwY5hchinDi6grJicBg81Op+1rcdsajfKpqpMDQEf7bWHmg3
YIwazGkslcpS+gfDzNaxbSdT4LK1Dj8909FT7wtAEQ2eZZD5IxM9CwzBPe2X7tj/9xrE9rJ/aGdD
m9Y4XzWVJMgkFN/3K0Aa5p7nAKlj89xF4ERHxK5ZFXDVSkVURPqkMri3/SUWVoxd0LRBiW7dRObx
8MYOv2M5x6nXYM7H9Ry4hMhs+bty5xPkZgf94IjB7ET5n9frZkdLuSXBZqBe89J9IvZSb4oHTsBs
ht7SjvA2aGAVBLcgQLtAXaHf4wbZG0BUIQqBueBUkkGLOnYguKz1PfIuF19A1WjJuktDwrntVaB1
rJBKubvRtM6Iu4XBEtVlvfEuEnmDgBZoCuswlV0wpz5pmfEO66Orp5lWVYYiOwBSg0bkFcRwl8ys
btzM3DoZkNQXHlS3w9cWceqrjpPElj8NgtT8wWWHZcd0npYUlxRN4dx5z71yPqGuh9ssFTbo0XYf
BvCTzZFoOSWPeNlekDtOl2b25mUqmDv2OqY9qo9penU/fjsmhGH0RAc4pCQ+rvhj5LTTzhTUIqme
X7hEBkIKMs2U9HLeB7bNCg7W3raHV24Nk6QD/UdUmirA+iM7cUW+hIiBWgaSaCcJVvmtrzfdXsJd
dOfzvndiEmv+AauttlIKAszBdKLCEZKOnxnKA674SySrGs0vg26rfm8grmyUcfOHgVYvPKTGhgUo
BEyJuof2/eKl/8AzF1kSpePd/Z4JsXRJUFLkt8hBowhuc88oYo4bqi41bMgJqfEUw7lpvo1Me0Nj
axAZxGfFL1qR/+95RGKdOn197Y+4R1s84s8gpJgXWtjmOkMI+kqyIfTkrd80TqHz/8CdrLuZeyRC
arnBWNAOAAIyep+L8Y6gHVOFKc2lrHel3od5UOCxt5a3vEcAU8nCtqSveDggI9mZZZlqXe/4FRzx
ydD8AwRtBDd1xaKM7lB/xPJ72DXMZ5BENA5QktN8UFE7fe4tAmc1zSHS5SkiBwa4b6nI/qUmtN5B
Ldr5rdBLQlhI5glfUpAS7ENRnNUjaFM0QaCbhq73XZYnP7gPC5x+iFSrVxNDUgJDQ5kEFCPa2R+e
eU8xX24xV2dfg4T3aSkA2E2imtj+wi8XeRCfVJsOXYQ81+LNehP8OZwtX/jH4AXNGhrgH9uPE1fW
IQVTTnE9OFptwZfGm8nEhHcvcuXMA3v4rgKhvUi6pHFPAIVupgoBYjCPx+Tvek+f8VVr5s0adCKO
6j12T9CN78PjcyXvz5btwqQxn6RBvjZCqSmr9FOUdxAvg8MzYU6jy15daOl08ZtYZECfThGeu9Cd
FMcQbYdtH1/vc/q8YSySJhe0hjQ/DsnezArRb2nWWClxLMu155ghjRmmWuICrgk14nHy5tgR3ybC
QgpZ+BxHwToOCGgKfE40ZBHR1fNvC7yoYXSZyURPz3ksMkMYBbYTo3UtFLBKZyurwvaE6vZM82vo
ITXpEhAaof+VZyW3uEbXnFu3OHdkpmOfxT47GHtPv+nJIGpYb2JDctNa6zr0ltLIE4UyIg6nm1hq
4HbN7F+Iwr/QOJ55zPhn2YtzrZMg6rGqk1hZeBwq4kpxxWTBjoDWbrjdXz5mZZA9qmSIKVT5lba+
Tk/y4Tw9a7TkBS5AIW/FLIoCFZ1QIYpPXJKWeE++euA501ruVtZ9xQH7vi18prMLaE/sqbkJ7+KS
OimdEN7JIJuo5WJIe8JSW31425KKO8UlJ2TdiJJTwpWvE61qIK3LurMqE+m2zIVsqNFMHQnQIYSc
jYZczdWo5ZXS0PM4IaK9NvLEUnzI0CelU6SJd4pb+7jAf+vOLgaFO0tM1IWfKX0tfqqz8pPSM6mY
KhK8pnigvxKUuU2OIgQSYm130TCaZVm4cyBtZ3Y4lznZFteSDMhIu6kGeCUJGe0iw7WaVUKQ5l3W
hM1Xl2T7POVQSOYEeFckZfvcVaM+qOB+99GYoDrKQgwnFsjaIWF9kUD84L9vMu7uL5waE7/Iqq9j
lJpbI09fGZQPuE+drrYljPGAKQAazPUTu3nyqpn7wyBPPAc45GEuGmfARtPy8iLKc6TDo6sGqzmI
3ERu5PqZNarBmq6vWpEFQ3tV3AKFoVge4LFWMv+8hBtxeXonvj1+7NMuiMmU4GPtIoUbWmRRTQHu
DTNpICwaCr7i+MPiJqUKcUzvR0HkueeoHxAftOvsrCymUMRz8QBPMsYDlKhGLR025/RTfnonrHm1
oEHUJp12YFy3i6/oRUDxbdmWr2xB18lahT0I8gBVkRVNEFElcu/JtgpY1wgfvCG+qt8vB7olqURD
69ajIBa8E5rRw2xGkl/PWQ+GSWa0R75udpXtT4WkZAWBU34DwYRE+cHq/VFdG+fVd2+GhjBI1WC6
2ecUnafKWWPPDEGxnOEEoYNXPQWjl0GBZlHceBfdWnPhBCJIqCzhz01j/TnaYH/dPhD8IKUYPN//
59giAk61+Yex4/kz+903Xv0NJ+o3P/OB3NdO7QS9oaTxFDQ2bEEy5nm9ksM3VPL5c5vbEVRvM01P
7bhAx/64HHLqs8fu7sslIOd8OSMjXHcnAAx+YgWTWz05z4tawM37IGOCukd4xc82Z/3TCaP98kHy
S+wgXCtpvyeeK3+4Ky72LL0oy0yJ7cDIr/vuFNKTbs2IwWGQSS44UnqeW2d/erMP+sf93pNyLykb
Ncf7e33uxmQRqMLnU2kEADfBfPHXAaomCx9dHbxdzhbNYGGZL3MQQzrq2/MfFnzy7QxvTFGNfkjJ
s1naCeV9sKqQXFgLVx0WZFM5+mvX09ZVDbnV+OQf0aTltHeZhU9177CYyZEGovjGsKaxdnGKK9Ov
uPfgnLJDI5tTlvym8djXSpSICb6IlIHYM+b60WtCM3mT4OvPn4c9JJQEO/yt6LFtHlqFplT5HcY/
+QreCVarNOdxnjKgGw9ULRhPu0ddpPlbHaeJBo3SESN+W8gR+jDIBjH0N9GSLwPfnxZR6D2k0eOL
bPwSGZbiKLfn+UOzuHxv93t2WvSb58b+EbcSkvnM6+JnKPJzW2nZLeG4hEmC0fOWkLzoE85cSoJ3
hv4r/keNVQSNSBdTnuKH/DNRFoourrwlpXpRWN0Clp5NUMStP+bcA3Ftuxm0/VU1GAsfqeFAJayh
9oQIQERfLPIG1i9fjPglc9LjBPFravMgkgb4ONmAo5yDbknfNxvoxnr9+5fOmfwrmoZFGL69DO/i
qwuF0ft9HJDhKaMLu9MnOSrFM6fJx7P+GOl6fuVoO5MsqnmXpf3HeiojPL7N/QuCuKdM+cav1Smj
O7IB3cyYzzqkZoOG0y5R9WwQu8fvEYzTnD+ipJULGwuBGI16GTexueZJdurHUI6D1Fo5fnHxpi5e
nzFWElJm1kwJitCSi60tXRB9wCY6YmCk9I82dSPUO6urwz3yBobEaOOETlwqswiSmd/qOrSUsLVz
d1qssqYdX1biK+2oGdnn8w5pPqDQCPsC/nIEodsK1TdyiEl4dbNvaORoJSSnQTsESQEk3y5Fpg1f
rkC/EAmlo940idfuUi5Q7aqQ7zFY2TJU5zWasew0WgelE8x8ucv+5Azk9raaOzaURVwXUGGnuZ3/
+SEU8/geU4T339bVNFAnDU95QlqAO4sSzt3z7tE0NbdVSnjO+dmoJfvkqg+jaPLvpB8rmXuKjhj3
d9kCuXaAlTmaGIzrK0SSJHHeWvMiaTzKt2alrWhDY8p5zZDO/rMZY4a2mGk5vJo1lgoAUPIx/eWy
kE8Ltw5n4w7ldv9+fdtMOeXQRNizmIFKp/mr8EhU/iJyY0LoclXQq0XvacQ/p7pNN1VuXFJhI9Ae
Rh13UHbutAJLM0mFy9Kn14uW2ArrsQWzrKDJKTKcJg3OH924MIGqpGpy2DeC5QJRUDQRGHN8uYaN
S5PuiknMIXDQNWd1qECFcs8nRRSwLXXvJUH8dDRqA1w6VJUCtk33jRwPDn0s2O5r+pV7snl2NG1x
A5ymuyyHSS59hryujpY+aUBamBwEE9ZrL+GHlDt3PjYyUk+R3bcG/s64W8eBOYgye5cnEJ6dV6K2
A4OUx/vU+V41uIoij8shLhV1zNUe/qg/vpyoTHKIl74+RToemYVYeRpGwOBAnB4vfyzGpNr9/bg/
LSV4ARafzrR39mRJVMVMnqI6XcOnj8A+Zc7W7r/ROgOvR2abxmxkD3ZKQiSVrOA8BVS0SvYNgpNT
uwbQsXU9QvbNHjlxFcexsTIN2rNVWVu3R7xaxQrQOo08wu9UWd1d7+iSP7FkGBFrjsaRLQ4Yms6Z
XVj0Rtcj/8bkLYW87DSzvgkz/+6HBx9B5+PUPlKbLEU0pznQmUpCYNXKJHK9nMYC04w4x2wCLdiD
4Oitx15BpUIGTYfTgPsVfbCDH2e+csbWRJDAdajh7OF+j0NIJ9hqY09tfk7PsW9tZ/h0j7hZDN+f
321IfPn5B322br5WHqxMeJkC+GGUgUKKFas3R8ePuZKsUSPk12wOv+eDvoN8qpa3zS6fDD/F//3T
+0NVOQ8khe2PL2BFyT67tqEskZyJ1n8RWr9cOkhQRJD6fC4/PacBcpyGpMyFACTDlUmwi3WayhnX
8IPwsu7BQWvPiIT3o0k2wH/U3d4vg9bnJLaytDHvm4JFKzMJg1GQqTPCHm1osjFidqiCmhsA1Fyr
a3b7iuKRhKIMRMFFCPX26hDVZC9qH/yii2+kxKaT5F9IKxq0YWe438ihXYF/xoF6a4LTYsg2QZe8
sLUMEk/hDP0v78tvgQyW6sretHzDrqiPH34YrBxMM1j8irEMyeDvsB++JoApr4MoUofCrE2ZLJ0a
97aglSicjibDbDvUe4HruJpwy8sfcg5pa1ZtzsAUwo+zW7KbVPxDyTQ+nEtrLhobrOwshgDAwWkU
yX0uR5/MRps3Gw/miQ9Z5hB8sK4e/+2Cx5wVuda4uyDioKWzK6Ce5dArCPjRnMNELw5PjCMMwg1Q
oiY4W/qoHoYYnnzkG7s=
`pragma protect end_protected

