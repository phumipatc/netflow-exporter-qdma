`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
W373UpbXC2jYVkKzJJkxjXwaqikiZBrnOqXXRtEXR60LVa0RoYvSA9+mfGgPLhWIjsk6/8nWY2MI
pw1lSaLhIO77Zp6ssLbzZvQG6SyejEhxnWrseeRn/9Xbkl8frCHSC85wnQLfAZCpTAbstlr80BPM
VT1UHwjE7MinTYvVTERkZ3tT0PSVaadKhEByiLGIdh7qW6c8qHWKWYNCAxBBZm4eM3DKoeyJ4lk8
PSYw+6xtWYh2Se7wbCifz4S3O2J/nO7XiLb6e6Ll+T+cfhlRuP/eD4nb/ik8KR/B6Hyr/4OYDQWa
JFCn9eeT7DOj4cebxoydO6JwxiRS0WWyBiHA/g==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
NtBl8z6dStOWc60Q0BORE83RGy7l8cpLVmVnLtN08SuqxR1kjlDIO2nrrGZ39Mq4jOyz6jsHCq7c
N7hLIg2Z5+xoeMJr9JvAdrDF4dR3CRK1IRDy0r2eQo2jhMNLFAhGykSuwp1xmP11uXyL3GRfhxzi
t9TbQtUqDdy7O8V5dpVKGamzvOk+FIO1UXQ5awvTqhz6YoZvoOIqmton+d2yjBZ7ce5TqgqXxj2U
Kwh8qp9E4wZIJj01lcuwowGa0+UjUbgw2cC0veZD+jMc3YH6ifUMms9mr3x4hPx2bzzgH6y3QEdX
MJLEx4DVPoehsuxl2i0tVIcK6dIAQT6yDElKGQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
q26riKejSoqwNyn/ZbQ1b1Veei/Rv6p05O6B5a2/rQV3SlPu6JOKmr6TSu7a3aQWgJ7/Kc9/R5VR
gUn3l1dM5g==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gVuP4XkTYeimmCwOseDRbc5IkZIWeTzCuIeXZ/F5Ld7359lwYK4cjb5MHffLMmu281vM8mxffrri
tUr+q/HNgk1CKfQEPwNKIp75O2m7MXePsLJX/JL0rpd/vHy3Yogn43KKV6MBzxKmlZ786vf3Mao6
v+jr7kKAODehtQfZGuy2LL3Qr5unu+grFvPkiRR8sZm1aUsY9wTAg/1nsWVYeb7sw1ru2rXHpnIf
WPC6ng4lU62/o0WThwYLyQMULVVES3OcUs2LVO8stEp7ems2dAUdLN4LBHJaAhFi05FdCz3t/ucN
3Y5CEuHhpDMfAR7+vuiOO+29QoJCKKaDCDCdVw==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
c+34bQalc6lN3dybyrjUZcFwOat8xFmddapGcsSm/D0Q62DYCSCC8ujn+YuQs/+t2qKD/M2in5PT
rMdsngCaWRrG835GbLT35F34q1pEvLajEH0nwRN2PQiMrVgETDmznXkdFbNNV/xBtsEl9Oz4qrVF
iHchKHsxmIDgp9IOSjIo2Fbw9IXaxfu6P8FT9d2LUqtBXpEKDol7RcIN7K1d4DfIVx6WZoW0kMNm
wIUNEBnIOjtqR7V30YSXoe2FPfsECV92u5oB93s8R/GaAY/6wWaRQOuTjnOoatlXnj+WINqkxI/b
hNIIHqcRu+OGakZj8ez0lY71sZR9si3pVnmvFw==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
K1DByxeti7W/NOhpMpHbDuFB/obBBcC21QtEDFnrNXoQtGMg3l528DM9W7ZTPlBLsoWv7b+M5ouJ
p7liycJzUKHx7uhm7+RPHUaWZEO060rxeq6i+n2N8qPlBYqoeVPi/m0NsT3rr9LHv8aqYuVkg3J/
teI+OG6x2ca0Rh6TmX8=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
FzC19Nxai/0dBDp3qWeQPqnYSPY+r8XXgHGgewKV7bwsYin3DoFZUNmVK7fzP/Nl0nRt4hp3o683
9dsGKAhpaVhrymE/lIx+jLJUBFy7Wpkmd+Lk8sUJc8+5h6ZGQWD36+whUqjnlm5cC/LA4p7Vxn/b
rMrrvydbFJRU5ZzFI78OfYshgoB0FSX9DRxFBvLW2orNxWTXIAkpX0MjJu3zdp7XFGFJrL3n5SQy
yD5c5fmbn5cUYhWTWuKv9Ek7McP6XwU+7ojLRFUM/7mmqLaE5gnmtGvT6I6IJ/MJFleeZZPOQBdr
sbPsSxnl/rUtCopS+xWPlb7I/cjZg6sb/gjaew==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OVNh6ox0Zw4yjzWT/GNj4Q8Z3vBi+dCBN+Psh+SiaF1Lw3dAFEa8kXw7xkuglDLMlQP9Vh5A7neV
r++abA+Yob9r3UmJZhNXgh1452JHh/c96UTvtqVVDD9yRo2Savt2TKKzFNYMCzlGGVVqgtrMMyo8
vf0gMxo3XQuA7p55bluCsoMkmjreKq7hJqaQCGbRsQJPdV5Fp4IMOsHI2PapjqiQA2Ze1Itr4lcz
tEl7S5P9Z3RLovUnvZHyef0S/UlCu6Fh58ZLqyPBkqkG10LL17PIpt4oMkHDa8RhaDdytP1gvVFx
bCEDKlHeAUDpKRqSJVFPxI4MfzY4wmczHDBitA==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
cYOzdjy6YkN6JcHdSTB0P75gz9iydS0ewsGgN0c6vpMUDquazoGCwk2tDlF5gmwBTWx6qJoSJvRu
pE6JO0eFNkFWy8qkR1TXaMRUS3X6j0WVpM0weaWmlYnoXNaoOFwlE34DMUd7BVad4slMWCLmTM6U
/t79AJBHcrpLH5HNCBQ=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
QNHAvwqamUsDs8pJkchHLNojBYJ4YsnB6D79z+zT88k6Gu7eI1vJx9tXIPhWV+GOTOK4lTPnaqw3
HEt81dOG8zow8+4PwUJs3gxAvCHuR7iHHPrv1EykB+HqZcnF14gXvmgjilczkhoArg0G8Lc8sdxi
0Qy6P7W8tgkH52xrQsW2emE37z5YCd0JzZxlVuLhpeAFcIZJwKEYesD75QGRHkcdhvhzhUHNZ3Us
RUZEU2H32xcvTgMhWId2mFXJbLcHcH3PgDFieYpNzOZHakF65glmxKiwunBfxe0Zfpi8FEDa7woP
J2TPuMgyqWBoXsVLl4P0qYnCh50r+h/qjpV+3Q==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8112)
`pragma protect data_block
97+C+KivMRD+P0nodJwnGLRqu0GAOmYiKvS6gbtHuXAvJN9QeEzW+kxtWtQHDWm6oOFkTXpiaIob
75U8F0TjS89h83xo3STZeQoUlqnXyPpyeBsjb82dJ4b5ur3SQNtMSmW65AGUEo9IfFXDMJU3zbR/
OesSNbJcwJ0+K6H8ZWudyxRUIgCD+Z8MF7X/OuE9lCjpDEpLtDii41KP7RQheFR9xCSYGp2WffOz
xvawlbFQyHxZXLWkiUdLd46e0H1amTj7s3rgUJ4M2y0Z8iSfqr2WlWh8ozACeMvKlyXiK5FuE06K
fuzSRyfXWnknfWO3+4B0XEWzMbka7p015J4o3SBu19Tf2hRz76R3u3XsdEiA0RHRFm5U951rlC7a
LV+JHk5ZHDu5b1VuiCMnY1SJGjPEqoySxkA3gRCwUjK3jl7mbuTpfYDoN4xbu3I3aXWLuCFhPam5
8QdYeBTu2WCs3uJ2BaE6sMI0KgqJZpZ3fBlm22gpGfjXDSggOJ4zTuOVp3eD8osu5fyScqjWJpsM
HojQic1O5Mmep0RoaNk6h0G6MP2KXb39xwBfoy31Jt4PEE5Fd3ZHPM7YAvVkYKLxIvhotDfd+eCp
fxWJ7Q/Wk7qGnu/rFFArZw0/mQ2vowiPtKPeWUezBFTyW3LuNBfGpGEAZXLudBh9tlVxzvBaXPdp
+aIaoek/MpTpwwv//PiV2LkKvlB+A5J7MQ/IFw70lf7U1DQE0NlKA3MzHmV6sukT57lkVooqu2Cw
sKLxv97s/4FZ7VpKrbYOGGvC08j+kNngt2V9huRgopHYmHyMxRwx5DDE7ClsTFuAozNzsL1L51wf
7ybj/f2t+EtW2R5DXNDpPMcpupX/UVgH5ZZm+Q7XkHv+GaIbXwh4iMid0Oi7YPRFacdpdLESgkND
LPRD/rfYO5oQSqCJaCerrnJIMz9jwx5jLSwMqXlXHMbOvemME4/uDK+nKV5HZW//4e44WTo1luIC
t4ZnT/5FAv2gebTgmBEaTXwc53/9Ak6Yz3pk35LKwSs9irFQxrh/qbn4+AkA28Jh3bqnEBoS3Uxe
XwTN+Ybhr1seDffNGeeO+HcWt8kfxXMA3iEp+RhVdHpV2QUUEWXxj+Vz6/8tC2G+dj6PexJvNeJH
MUEOdJrH77Q4ZGYw3YRR7h6APH4NzxyCKT5DxjO+Ybr5zKckfkr0Jvt3CoKpnQeiiX3q5cuFiRCL
6AMpLZa/bOxhj/2fK6IezSaHZIe3DXSFen6X4G3PgWsf2GEHcZSmDxXV+uT34EhhTLI8DyBnlrkW
WoSkWpiTSHAdUwFTQSo8/UeNA2GrOLwnhoMps4P/4Hh8dOAPfh/LqX/YpiyDi7R/fZkQVrzxNs+w
UYUKfIaTkwyZQoHt6cf3rRL8/BkjV7+c7uH97ofGCb0V9yTSXqI6xdH0eEE0bOyu6wwdwxE8l0FS
w6EwaI7JMBuElL1W3myHfBRn3ZUKv37/eORzyV0wVEU8OkC8nYJ1Azn4kWFJ0REotICW4v0Z1Nz3
WsAlE032DWcu9x9lM2h3f8AzCXX7HD3BMg5HPdmWpapD4DmfPE898DtaTNQQvM2Fn4cVEvJfr+r3
K/ShSq48PTO/r1JX1l713EhykCuDQi0w7bY1UmA3VyRrdflqED78jsXficJFEYnGVicmgnf9GlMG
QUW+51E9OlF0NIclkGJ4tYb6hOJFdXdgkS879qQ964ggeX9MM/lY9w+d9euMh3yKzbbTwHJvTQNb
ar6nCVo9lr2gXc5awsergTMTqc1HhgKyOLSJtvJe5RYURgHoFpTHNl00Etw6V2aDgoGv4f/Zqmhu
Jw6U8LOyxnWhDQGaYWRlE2lzZXq9VkATrszY16FKNvmxaTFg7Yx16PZn1C6/Jc/fLIIXbmMFZjuO
ulYt1NXVZQXZ+cmUWQJ8dM91WDvAVPj35AtCvXOU9fhdC4MKRcC+8pSDkUvmnxt2VYg1fYlg77CD
/DRt7mHmb1qIEghbp/EYxH394/S0MDNHnSfccHKF4C4W+6Mpwc4JTuAiCX74ZolLrrVltx01/XGp
0GHqGVpTzNSmY9TSFhP/HUmKMdfUVsnDX7S1XlD7GWZrjiw6q/IPeqbEG3hHpF8DfLXfeiQV7vvy
YIPrDcL//6SAPHREBEtpH7pyjCeMUu806fXOmgnjuwRCQEP++32w/zEQISgfjcWJaIIgplGy/34u
x9wMtNPlukW3s1hy8Rvm1mQFc+pBiLY1iOO/zByrwY8/K2mYMbGkBv9Ajt/XKYtG6vqhb9/hAQo1
rjvtG4pL6dqNQebC6WFZAD6UhRHM5nhrg24KxHPlvORroCj90wrTV56f24v4co6meNImah8a0st9
JMCHRqAGzaLE8bMWRM26D532ok0gV0g8aayqP9wAi/E8FYBCCYlfNPQaQsjhlny/++vuDhCMOWeH
w4+5r9raH2sw3V9tP5NB0sP9UlyX8SZDOdHLeZDnAvbU2Q/04TrVWNhDgkqZwgHPI1uSj8dVQnWg
5MYd2eV+GZXdQyMphf8LsLyGRAIAqCVV+0c+t6LDlEat5dLryr/fP6lvk2QrRwIzJ5JhkEm8q9Y+
11+ftTJ7AVwYK2TuIJroIm2ZNgW5qpXwdsPJTyHQZAxIYG7AHbs4heUq+3yKQpXEEbbVAXM1PpT4
/OHKgXiinWM+ozz8Embb+rTQNT3z63pWu9ues95OTlXs+0cu0Q62rUYzHznUJKGqlHHpx5eHdHEt
3BwfEOfwWT0PtMrHJMP7O+tGm8BvijZbbA4WVSiTa8EakGl9vHbcpqMPe/vkRpwg1VPqlvveA0rc
y7/RxqHMyZPIhjbZ+wTwxaVbDk8z2nM+vIAFz/IKZNEIJpLpCaUZrMkw9uVltuDOS+yKKg52bA9w
ZMN6Ghz4VbawjmlnUdKcO8mAAaI96zNS4dOhphaHCqsanIwuQaGImW7WRynHmPch9Q8IpN+pAux1
NaolrgqbBeLPlzOYveDUMNwBr1bdsijnF7fUZh6apDJBskBtIqNrFlqxXG1jzUHp8K9upnfsF7Ev
9TsLZb5uPKxLM5GvpqxUQAF+CAYPjPatGsMZefnNZ0+EMETGipDohxX1AbGTwfDWsutB3Lt60HFa
CinpeeynuLehO4zlV4NTthhFBNg3nd2QfGtVEnVilICLZ87oXhrkJn3W43vH5f/gxkPSHhwAiJQ4
MtYxewOCuffWLFhzrN7puVdXoDKdjx+M24i6EdIEbZeGJWlDU8Wj2EUfgfx/7Ia8w44uDfgixuBf
P8/rl2RU9VN2jqkLBw4Cer7G9eGxN/LMrwUDWLqgOU12w39TKyCf6uUGjxou3k0TWNeBN8YVT8tB
B9Q1XPtpE/0iwJ42rH04EKscRG2++pjJaePH76MaT4YgHTq0RE3TpfgZQCtg95vFuyyGYJPBKGjk
k8Md1z0XP5ib1humGj0vWzfSpvnrcJGRGVPkd9eyX6SQoAFpplSDJ7ATk5YbpW+CwSqA3zvKpyMN
qZUfehX9/QoFcRw4r+A+6c5wLZoW8WlI7x3NCjF4DLLTzdvqYLxvywd12t6/bHxj8kZVE8wfdsV0
ehIi2kPnGBqza2NjRx/An/anuQsMFa4BSBzjy6hTolw4ghKhmGSMf8Wyy8RwLfV5wd+HSpH3S/NA
g/DIbV6teeqOiGWWixgcskq+ge/J9MZ6+eynxyQWfw7Q+DN5g5siBGZGFum7CzTLB/U0fvgYFpfL
iFb1/mstBr/lBdb5rkC+9is21KBrSM6ys0Z5cBm9JGk2ZyFA76haq9mc4+FDUx+lhlFNtG0gDZVO
6OUl0g8FzPDb2DByBHcxpyVsw55fvFYKl4OVSJi3NX8a/uFE0Y/Piw6vLVO+SIOM1gBibER8NRL1
6uU8yrkCjE3VmIKmnnVcl8YH6kkFzmOZtyj1/279NOKz64Yvlaobsy78rvWoKaLUalUSCH2qQw/r
g7MfQP3M+rACnHxYYstfu4SmUp+wn/a2GEZy0E9vSCW9kKS36ga4ECrzm1Y39HIUj43FW28Dau7L
XlurrNV9YM+dDtLS4tgcP1e4VQ9gwvX8cQ4oCJ2JU6/2lrQXl0wGcC3n71bTGJy4vqsORrwLgytL
6vKTiCt88bF7zyObFm5ciYKYm5X38IGjH1MII9fPaFNtCEX38ZbiiD9DEFeVm1v6wkYanlybg4bV
ucCK772PmQs4I9qlJXpFjX4a+xLx4VHbtbSJ4U3XllleH4zcxezLJRDOmEgRz1JFJ9S78So1wdOU
FIAXSZqaxqc+i7QpLTfa5fzYcPTGuDdZao1qMyKVzi8UGaRtusVB8vJisbLqxe25PMbExcZP/ULB
VJ7xTfau5ipa2eAxYsOYNweDL++zEauz3gpDZvmu8GgAPc8dEr3H0N4WkyYl4d3Q6gvYtV3BJ61H
kt4UQ0veA6F1yNfr7LBGII2hcjQ2iOX1uAGSzyeCu/zplUASz3NYK0QrCFqKAF/iYiTr+9TJybE8
/rcIowqStU4RIGTMwM3Wxq+48NmzSF2ldq4EjadPG0IsmcX0/5dOUvKXHUgS1yxRRYhshvqoUHh9
JM/MhKwZFS6zXMQH4MLhDYRxgrUphUpueD/VEPx367DGyDwR3PIu3DOBPk7QXNzTZY699BsmkYim
S67ELCyRpDbk6jvMP3SX5AS8C5EABSiLwmqIxCznPZ47uJSacc01mB+ly+6rF3Bqiq7bjqMKqPCD
gHxzsdNot22zNCNymx/WIePYMht9Syas52K/IzwALjiJn0XCkmZAWpmuAkGqqR7c1nGsHcyirrwD
ntfJgiqLL9HJxC9hbo+zrCB2kUACgpE5VhsvB+cmT3rG9mOhd7aKMZ//eXzMrZfv9S/KESuB7BvI
8LA3kLuaEKMHuIopYxgEPle++5RvXu+suwD2vgvCNXztj4v5QUywfMvog44+gqv7FPStn6EXHwBW
cOgYPJTbq2IDuMHCZLi6GS4Nstc2m9uLfJ1isT00u0OXgPOkEfVooIPIITAw1XHYFY50r7/qVmwO
K0uvPBzRNBCETPrhtsUsfXmMvmJuFCGoS/bGtFk5h0cEChsPTK5ljBDrOdWXZAkQpQpPvi7KvYB7
nXWqz2GuQ73s96ZMI07E7M6ol1WAMRHPNp2AoY+2v7ICEvGAFur1EFpKtJeq2jwIvwm1sQsxF9TU
IPc8VMzE/D5sMTWp+nOhGUSVt0HT1EedHIwzKl9Lefe9HCeOju4P6NSQdCiP+pmR5JgDL6Rdpk1J
kO7JZNxY3M9Mgk1v0i3GOi4k8mSUobv9K5GWdpSiyt+wxDu9O93VCwCwosGF7UCJbNXZPOqNcpLS
8n4e92ajx11UjGAJSzKnZe7xOSmadWruDxSHg3LxuPswdHTmJkTAZySnBMcFLg/IHZ3qsf+LP+8t
aOtOs74pFlPfw2Ik0olS1mEYr4YXkHZijLgTaNTJKLBSvIqD4eO+BdZQlrs/x1DqvqVeAsH1BQzm
g+Aw+CD0caj02G+e7gFdxaHmwfydGT28OnGZBxCnqVit8ahmajW/McPeVsVmV3e735l4fOzsRaUG
VoeDJwmODpzC5ANoH6rIRp88XkPL1FDlEZCe2Cl0wkw5n4aEKyWAbThypPmSOU+aWqiK79WhXE8q
Ztls484MqTefy6DqBsjmXRvudzvUK3nU99fwRCz3CJYa2yNTTPmBTOFiDnRUIBBQcPDGx37QVHUE
x+QRT5VovRVwuh5wT9tFYgN3Lnz9tD+inhMsyk31sZ/YNjerYhSCDbZ56GRvxTiQoQxPOUF8TmY7
FZNr1NK+924JwzuDIePeVy1MXkJlEdWuPvxuib6snTbEZT02p5hMBC9Vk8jpLzr9w/amzLk8E74j
E9qejS8u3Wt66tNrCeGapcZsE0yfVuTLEgh8oOsmhThtdlMJO7SytuHQbCKJKcQKA3TLc3g92VFh
nfliNEXH+D2oZXoQADW7PqxK9taea+2UHS9eVpJoX+RQAQk2FPZMX+XbVovAFnB6NPkg0WZxNRwq
pcUVhxazP3W5dVCRsLHPWCuPGqM++kR1n5YriWgjw3+Z/y39TVoCMZA3juV7Ikx8vq2GxJfNdk7h
bX/3lEVSZLm//ExHIP+AnuK7bfCSNd4Dc7eyCjdG9/W+WomcGx4SmHuWaF4Pf3QfKQxuVuX7rt9t
IH6ApFox8nLHSSX8quRyqZbc6+Q9nF3/w5RrADiSwOQmTOwaDfMQDOj7IiKT2DNetyZ4CZqtTVD4
kvDEgtOdBOtpltw1Qrsdu48yaxO0QbMFzhplwbCtTuK7yIAZJGbzaYSaPHGaMUveM2LhQxwStHlp
ejw7zWRkH5r+gfWzQ/4oKmEXlLaGywETEn/MNhEQnzka6FnO9uKbaqX4qU6g1yvncwlQH6QqUrU3
tAMisuWExsnKyopJZhMX2oDqVwIbaZdwze8/3d6NGnO+WUY5Hne4d4/MZYGN017U6Tzto8ZSAUiV
tp0L6XDxdGLGzgyq5HC4fX4eS6H++gDqb8CsL4lmK3MgRbNG0MH6AhcITs+YaxK03qeRPkhFPYDy
MMTiwRmlUQ9m9BnUz4HQ0CcTFYEjJpMn1feNJK7r5NYOndH2aclFS7yhai8dKZjrmP4HJ4wb72Bi
js5+grSSd9H7eAz2CuOxtgFv4DHr3BT8Op/B0jEHiC7LMlefRvzt5ldOpJoWYk/miaB118J2GQ0Z
rOAezWVJYA4iaMjgKsTtPq+lf7ax1g8Kv0ASikwNmAHHOyDhiWSJfGGSPI3+Iu7gqMrrhqJdad2j
wWVtwQdL+C5rRhCZfuJhvsziqEx9socDHonbmOZkUBU6CgQf2S0AtnzTNSsA3U++PVudePXr5Iac
kfQ2BSQ4NaqiYbppPPVV4ETAw6MSFwTYb6wh0LyHWHleQcJTWmFpLrmGkQmsBff0WkNkYbbgsXes
v0UWVs4rEmVOzBhPr9SjtVccBCQjxk1UQ1qL4h22siDuJM4j8nzMmP8igG5inz1BwaP6WSgmqy6V
8vUiMjMfibJsGdidDoUs/fbBrXhni6HH1sU5unPEMd4ENTJF0I18qTcYiox/4+ewQ7YHTzwTy2i8
xT6nyMzigZUc+PUi3rHmhJd1L5BcKX0AICOppEiYt/nbHjiddncRUqI4WxeETpK/7NdRpZH7sqcI
73ka6wivDgIK6fcoymuMX+7gDrMQ1pK+gtPMtWiFKDBzTZAprDSLqpPtmLtHIssj2yw9xXqm8RYH
coiF4LvA2Ae//p1+a0URqptT6Sjn2Ymd5PTx+2uI1HapajMrIMPSN4OzaL3DPEVupG9j9U4QrnXr
PWIkW5dCaaszZlZzH54rBrtDEzxs/hZCeeGKIeP92ZWNKOrrZ7wPDFLT45wfUIG93XkR1xmmyrh5
/dV1+N4X6Hmg4E+G/WSpdg+ZyTHY/w5wbmrrwUXAbpHVFHKVXRyVEao6QmEp7fabL4vGXVMepfwY
CXLqfmqoSZolPG/yxjU8vTjCmtgUy9+sgvrRJVyS82vmkwmdFrXAbQcmALJRlN5HNUqXXbb6z3vX
n9l5RorLJuc+wxesWQHK5D28j42Q5eneu/DY9iKh7vlKT3WDz8CCXs8aO/74tb1WAl17oXnufKwI
clI9WM1BevSAyCNSt/uO7N+cXDx9Q5IG8+v4OXXQDVimPM1xBehrx1OAQvuWir/rB3+E7mKlbu+m
Bv9BXcnnFOIyAQE5ZMOCNWmozqXE/D1t0X0Ua2s0pznvxVyP1PtXpkIj58BOCl3yBg5j/SOCD0ij
gOGQPG6OFcjv5WXUEr4hNSu7kEw0lEAIM4owoa1FT5aXBAOwvVn6Pa5Z1wlXPYxJQCXCL6gDmbrv
fnk/q58tTXQRpf6UvF6XDIMfm/BqroSndeyAX4cdwdR3WNdgCJ4MKnQ7DtK2KtSMUe79JaSbYdNj
NpgXW4POqeQBwIVd5vTA5O22icdOulM3rJvNGOMWYHaA0n7ZCojDvtYGSupjP7OJONYFhvmK5GYx
cXWkqbnSOUrsfQQX0XJVDXmAX0d3YhewAU5oJoFyXgZA1hGCvLFKJv6m05QB+6hXI1771+Z/S5UE
FCK7iXR4l+wQRICUfTS9hSCl9E9SXASvwXupi5G69auOBIshoeNBllvTaQ20eeMs9xqbWKd+qliN
IGDYS67B6XYFw7mH0lV3jV2A+8A9fUBP2MHeB9+F4FCFuvpAZwLSkV290Y8rHyg+jYX8wTZvcaIT
kVZsMseufyPIY09p9h6piXRdA2UzcM5oN3cgVDVarI53dOII+ies9KhQJZdJk+r6s41rBL6aei8O
zMvwi1HSBgFMabc9V1Y5KaXYpxXzJlqnmtVaxA0t3aS47LkEcoXM4L9p9VBnMW6AUCF/pYnDcQlZ
VF1lYY7hvmLrCZ85P0MKQBdQuncZUKKJl3c/ocfukxUhGkZ1kGd5RKI9CtuABzGJq210DJLe1fj0
ijSQauLjdgsG1vYnHDLDe6nhlBv0tltlnYzTG1BHCvdAvWZdD1b2RCTxd82tV64YJa4Rqc5F16AS
9JblK+g3pvu1eYE+X8KWHyoEPxZd5MaElpHg08QFu/xCqWS1dBYBzY/nZy2P3lQMeahF7OkWmmk0
swyiaSnbEElA3rakzjDDHrTQLlaU6X3B2LViiIJfB6KETl6kpSAldSFGAwrxOVLoP3evMpy504EM
RnaXuDpLaiTVEHEdb7FXFrcv0nEKjkPQFo0XlBpYGXwbHo0zzrFuo/vZABMXn4JkFpoA5odlsoSW
hV4SKRkouMTGZtWAq4CbmCetQ5EhqW7l5A0hqRQkYGEdcvPx+mtqfKWig2QPbQ5REqrOD5emAoDN
3dqlufw9B3eQY2mCLB8iJUiPThtNwt2otGhz84O7ULuSjPLqCugHkL12qJ1248/XZZRTlJG2vWDO
kwlidwfE+vAZcM6p//V0ZWd2AnUCHjENakOu6IOH1lVuptGrqn9zlWw3OwAr5XRabnQU6zx2oFtI
iJHoHM9GNQRmgNVg4hrOq6u9Tc6/t9xbs5ydQHl3nwne4WEMqP2tH9Ls5cf3T0LupUb+ROyucbSj
S37A8bZpLMFHus43fSQ6l+l/VrrkkzxMnVCbEGLED6+yIpC21DXmyT1L2B5TyS0w9GcIDHCkzgJr
DSIGN/JADMZDv3rcEeh1mocIebEmVQqbFWuPFzj5ofGPgrTNfHmBNUxODy9mmx3ZBd/3AuqLCBBs
8UomoZjgMNUMd6Yw8sh9ntx6Jd0c1PHnZPnhdfzcGH/BFG/a28ktA4jgUbN4KZSuCem/zBv1TGtk
ohWVLT+VBPgzrpbTIk7nh+Z+8PGFTpctsIQNXJ3QZ977JK82Hh5KE286IuTsCsb0CZZurl4jcHSs
gLxE8OTapHQ5BcBsFpvIJO6G08HSQvxZuhh/gz01V1u1suEoKVd0FOGH2k+68YCncp3M8OTgN9Oe
T/zMgTZD7ggjKgrqagMLSQeI8qeF1YidMtgYt1bnJylG5t4VaaFzWywai235bzKGMxp52lUjbW4S
NmLeyR+KyVbUaUprDgfzgJOxSptaN5LZVLYXVw+GoML8SfSx6WBbLkDxhVEweOmNH1HB4ig97HDa
DQ0bAEShoCzw2GE5p2LpzpBLdIhcJNi3mrcNtKiBHQbuJRLHUf9hlOZs4ZughP2jxdUfkZrwJ7sa
uSs+VDN9nMrZzkFAssrSodsCSr3j/NxJ6TsE5vfQh0i4m+DfuOxZJV1kzRNNPEV1vF2wouGsawW/
jTgWT1fS5QW1YZP8gP66Ovn5Fs8vC2aE4EGZgz9k2nqKyNBhHaJzUqltdcSGKzrBzqFHXnC3OCRF
gDXvQ6wcJd307l9oZFR+sqZ3nhQ/TbeDJfe68vbzpGTI8z9XH86P5NX4gBSOD0mTa6mVHnT/R9Fw
9m8PNDrN65d6ENgJmxKnCNh9191TZ5hb44AdasKvcl+84E087+V0M7BqV0XhwyVHkJYUhhHYZ5Zs
EIZs+NPCIzRzIkN69eg8+Eh6Ko1XL7QdPXShep7bryMWXMAD3iZavuEEEGUJUd0qwAG7BqAJcZLx
aylq+Z48RPDDaxQq/lRLwmR5VZSEGeS63yyewYdgb8VXwBtM/poxynbI/9cJgZrgcL4YzIcUpC9d
HDT5AcNkT+SEVQ4qjGeTp8Io8Y6f5JccGm5pbCbVoSSXn+UPqiVWdd5rkCkKU2IoEYTyz8xzYNkF
VLDcg4FAPCwZzQ/okwt7AzuQND8E1I8rgjGWQX4MXdTGYl+E48jrz0ch1G2lYRtUtS5iA4zU2r1+
Do2lBBaXb/f1CpGzKFjfgU/KVAwGp7/LhEiIsjINfRHUPwcFkEiKCAV3lnz5K8hHkNn2Q4cDGSd6
cfq3ReWcTdi9mrI90NGiPogRC/LV2kOjT1i+IayUKfkqCULjjkG2Uhv1oia3nC8f0X/m1/z544A+
1oKutpJYhEtCzKH6rvyxR8zpeX13Ac7kBTehe7I5NvZ6Rh0akQi1X5UrGycJkgam3rDuJLnzJSe1
EE6CHUoIb/9u9qczubp5mm6gjzGHfuTjsxa8J9w1n4qAtdayhjKpo3kfjHFUReFJryS6l/dXJhsg
R0VvzL0zoXyOuLCxWxyDjM7LlIYe+kl4RO6J7tEVwax6l5q5xG5SM+t9NOzzmUut7PSymN8uGb84
COgxAiJ+421CGUQHN6Ucjs5Ctz+KmECc3M+N+jILtmDbJviFCxEHoJP9u4m2zCsxY9o0MhMZXKT0
wN0oF00sj1loL0N1dlPHEJ8Q/hriU2yGlAXw547boufBtDFKpK+FeQyFLD8LHWOSW7utQ3POz6+Q
QlnvoENIiyw0zibzeHWxEado
`pragma protect end_protected

