`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eP2XARyECtfz4gVpNHBXO1U1tBKeVTpIyNZyPnejABv91raCYW/I7Vv/uW4F/lcVuu3SVMyVVjoE
ACLcqnaQUoeHKUUAAjv4LlyCPJHc0TUvdHsVLWHlNpU+f9ZdtXbzKCpKSPmJ49rX8y9GeVLLuJot
ETCV2BSLQFy0uGaoV1v581lWAo0FpAzytpdHoVkmL8Rzr6FnSnHe0BJKCe8y+qmccMtCm6u4QD7d
L+hZGdI+cT9Tnsh7B+f+N6eMF9gHM6kTNGlrfCyzUW4gKIiYcXwp7LcbIsSvto9mNlpt8f0RPokY
giPK5lp5t8GVLC5e9FtmRDmfjHv15MjOiRKq/w==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
ut9xm7d3VCJIbm/qLqpKdUnbBi9nwrCpf/xSM+Bl64Vp+Usj5lkVcI9O9GmxCaPSXPkvmxidqWID
ZiyAxtDr3w5BRW7nSjXigQLLnU6WlOYKmUkmJBgSpjVf3IJ9jM6wqRgKg6f1uIuoMwx5gzJUHmBb
VO1bxqsPqhl3GjjFI3gctkAVKLzZronRkv98VO/iobxeRGBQNtnwt6SRKwzZuXr+fN7pIdGVYXW3
1l/SwjsT+r0QfgHd6cJ8HCFbevlv+YiKpZBJsDlpO7RWDr/dmFOUkk8mx3DuoDP2xk/hfFo1TjuW
XWAjan0m8fd/BcCx9kEbqQB4sYNFRKZJrOwSSQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
apYonoNAYkxXZ0Pt/NU4bfuHAUIQ/NprFWqqDarsclcXjvikBTN1gZXciLi3JNlCquOwQHMfAxkb
v34pQWeH5Q==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
fKEAsC3dJCct9SPg0YqUm6J83ZOgWm3lb94nV7AlVytnjDWs/AuFSKdxtdcIZxHmwNulYNJ5zcUJ
9dJe18DnXZ7QH2LoGeJRBJSAn+nBfGTgZlxIGAVL9GCfKalZiC8I46Lfr0kE6fPmFcuWaoD4SYTi
Ewz0ohfnNvXPjPh0ODly3YJoRPbjYReNGGbNoNs3plvDOQ/4FgrrI6qpIh68lPZX2NEbyEhmfRjd
dXlxjBlLhdLbjKFQLi0hLZmAeFuTGATlQ2AYbHLuhYBrBdfAf2+/DWFu9P+CflhLOneOX8VBZc2o
IWGH0SlwCTpAhNSCw+5yCYYA5sB1BtZB/OX21Q==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J2r6M9jNo+BKj0uYcu1hKVdfnQwACgr16QUR/G4eZ+YsJ9IdPA1n1gpqC4ahhJfQO3TNBHTVHgIA
8RPZfcpS4pyNzqPl/nHT5fA+rgwpqrGqHgf7F4ptOFJfowyFrptEJKolzBr7DN6IGqGki5OLxrDW
9Vt30UW2e5kmtGlmdm7yGlu52tc5OhdCIEUpAAeBhSoP4697muvEUC3aPlReut+uiRRL61GYahJG
X2TT/RSyTekQcA8Ngpgh2Tfn/CoTwUyyn1OuBfiPf0va87WELb62p35fooK3FQdajaNCXs6DW9l7
h+QHT94J1sGpYUnlOYKGSkKK+4mY2EPuTMn2Og==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Cbpg6V4qNmVbBV+sxbZLckTTRHtYvenm4c/up7nxxfseEI8AZbMTEokBx17bt/VClZfQmTZvj4r7
LMl+HzPklPwL+Y9f6iyfDoZ9gKibuYT38n/bRw6smxVth568XvC+oaeebU3SJdvubBJFNAe7eNqo
mNsF3e8BFQo+aQV+6kE=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
c4kRcmN2aDAcLaU7QDgSj/bbeU4zhClhi1mQbzFoCmzZ0G5y2OEaE+zVlo79d785lnDlSr95Rh0d
qqXnvSCYh9iA21ciH8caW6tgNGlUXCMzn4B0Dl4AXF2RsmgwDb9PSCC7opCEZZTpif9SSE2AhYSl
TuD/ctANwNZbpZXPcEL9m2JyKAcSE5yDbSqG5umWPIlq6nUIhkq0QPy27GXtOVFFcOBg4scurofz
Xrf97U9X3xBVP+FdwiPS1uQW+EY1Dkdj9GOJJkwOaG1XZvcKnAReba/mVyPgLQ4ZOF2lHciuERwW
RO5vXVVu3uSTqAv3OkBMmNmDs0DQt34AfrBA/A==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jHyIoO/6QVLoDMCYnPKdtXRd2Y7CFU+4dAlQ0x3vrVYMVKDYS81KKtN5jDHHFFMz9xfOHJhtqcNz
oMJ/8EOBrASLuFiM3Hlkl0EFa/UR1ClwrKIacc9VgT3Qdq3TRpWCcvoGDeDJGusPLYxjioApJK+5
1tD0NqcB7ynbbzjAQQBNxYAcJnWj/tOHJ3b6iB6u4YwGWzI7kg5d7OH+7L4+e/U9X33uHaWkJCHz
n9us1YvR3kwFb1rlQJVi0zBeLfy7CeG/yDK+eygL0C6vZH3ZI75F0Gp/kuu6EZF7jvWpZ0dOPkHM
elpdVWPGk7LEmfR8vQKecrudX7w9xDnkXhEgqw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
lbkVFZGOXfqgkW4N+89mwYWLa2WX5NOA6bFSOy4Gg9+OHALBTmQ11ffJNLqr4NQMiT6VyunixpOX
H10Ayd8MAelbAMke2bLJ7ZCUx7upSP6t7+/xMAGYkD722IyqVnXdQk4Hj72WLjWR/WhEBUUdhAFZ
dQp5O+dO2V+FZHaFq1A=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mx7Jey20IslX++MCeSlfG5GGvG6Xa62cRkfxHE8wuqYRgilytj8hbum4X6zBYkzFKr9roP9idLOq
5rXszEsx5qpSV8jtHCrakRvcBXQDuzcByBV60dBusEPTMYxxB/p93FzzcyuzCkP5to7ZXPC7JkXO
fiyomRae+pWR9tG7xO6n9C3p+cieB7flrWEeNvlkCfXDYzWFM6vIjyhMFJnsPmdZfTtJhacCMi0W
RMtymeCrpUc5h9pukzVUjfIW1Q3goiiAp0BmSLEFdFPIsxtmvpvzuwTBuMEfDite5VD599VRpVj5
SSf4Uy30Y+lFaLZYcthcrl3lX6MugHjQfokSDw==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15008)
`pragma protect data_block
7V9y384yvzGU30MSZV5o6e7in6QC0r5jpOr+DUjbBMIg0tu6ZW2oGm2qdjZak5cxt25ElGd22dnp
M0vKyjKMrFrqDXG3mttWWvtM9PSo+2UmvJZzzDitDeNsieyPECdm7jnrNfaWiR7LwXQeC7+L6mlM
UyyomZPlRbfee5Adk4e5edK6nYtgsUNxwgRDpRQN67IcJ68i60++S3eE0Z0AHOx6zpiZ+19L17Tr
SC6/W9hOJ2xPaxomgRz6CR4a8LKhOFjR3esgr9IwZ+XWDws2s28zH/bLVstKQvVnwZEmdC4cpYVP
VMqeOVdnrm8KCCvUQD1EaQTElBfc62MFdun6s5Ds9f+nyE/02svqYbOHpAQrnWEYzoMCa/1aSEXj
zqj8sYfA93OGmzpZ1WhMD/8Iacge0MXPXVnumYsKOShC3a6Pyu/sPPOfglrn66vid7wnOm+SIVBn
Cj37Lx7N9R8hXxTxsCFAj62pXe9nnSIAoX6p93nT12Jq5TY+jIdtQ7xEJCSDWaOoLyuIAqKN1kQ0
qpRXs6NmTDBiMLI0W0DVOIRAjPtoqfu8XtFNOdBi9ka5zwLnlUr9nVVuWkVhLNGUOBiXqYyHtCWX
6gE3ck8i4L5RYSyErYCw8AZKETc5/q7UMceqQb3pX7JHTkmcG0tdvLbuP+CPAWNfBBpsX2z1uCwi
2p21HdQybGmvQB0GPmRzMYD5BCYWNBLpfspgcJ6jj3GQpCzi5zdKx1w2B+F6hvgtoYS7bzPgmd4H
ylyU4sAg5YaCKOPeb5eGPCCAi5IxayPVEKAetl/N6XqqXLCdRUL/dvdmKbDUK/kJDc85hWUu9bG3
J1eKOFuQo4nwQC5bSM+Zlm2GQCn2oG0hCy8EboVO3/MS29KBVX2nlEduVJBrk0thltHg6tqI1DSS
RpA8H/rv2dCZvRqQVLsWdU4NtZPORXDVTpvx0mPKUkdsGctxbDN3fCDUC2Yw+9xV7u/KMcO4LUnf
vFDWuKAaZXjtOKXzEO5cyUpg/Sedj9KE6qUtxQCbIYKR9YNIttFYGQzJHDCmj8jXOL4h2LmmfM7Z
5GQBQ7qYAKjxsOS9DPb2o96JBEqKrAbkf5CY9ZEH7dCIiMvWFRLFwmCfhqqVIodabY3mjdhEj2UE
zik6p8b9EWz7eeQ9fjCLmdP916bR6i0K5T454IQtfn0Pt9PI6K81jy8bDZ1euHJ8Z4+aeM67Zp7c
y9745qc7kyVis+bS8sh9zZTPcunOk55VeSCmYjHCQWdM4YsghyPdt2yUcGTKqAAZqbJ98oPvX25R
D/K7BjMmxfdLEyseu12mO4PR8DR581JApQA88nwEZYQq+QcyR+CshY+GF3jYTYrnheG+f72AxD4n
8kYTMUPSFuTdoEGGXOes1tmURR7Cuz+0NF9kUhDVrKWs4IIgg7td35BJpDUa9LXjewilCRuR/tDv
tgG8tWI8Jv93oPrf7aA6FS0QFGrWivXw9VFxVwXYKuCwjN4D+u4I5SrxJQij30fVFbwIsT7RlHtu
tq11WpoestvukcuiM4bo4Q2Csnwefcr3d+LThJlDg44piDCKU1p+2uvM4CkFtftUG+NL6S9SM6OA
qFAu9c9wL9MgrTM11yId9IFaIsdhBFTUmyT335RQr4qyoywRd2cS8VCTfhM4YMpx+NnXbOXH5J2u
iDtZB18izKEm/AbOEJKnt/bsRbvhYxL/GWlMdHePXrjDslNOTbv4ZPyR/7UdJE6SEh8RoKHNfHJz
PgWfeytYv4qa2Pdoc9x/Emw2ZctVzO5UFT5yaY3iAVoY4luwQfJL31F5at7QEKYaLwwsH8quXO7c
EYo708ENSrbRivKnUpHOD52K/85eL0JFlCZptOS4QxGab7FWAxxPKI9GUKPgwvQKMSxnsxQ8yH/i
FC+zB2z311Oqh+miy8xHYSfAM10vf9gW4WCbEuFEb8AeH2g9cxgwaCuBmOREQ0Hne4D32BnSa3sQ
KaWcV6fZ18n8DsVtOaKW2BLp+G21+UxyJV1HsQyP8tW8VRxm9bsmHG09nQaHc8WfxvnOO6BG3ZHo
AlFAh+YOD7Cqrl1ZG1lGAY3d3pcK0dNduSkZYcxL3cnUFqksl8s6LslE8G/HThDaer07XxXxSGc8
g4uM3E1W++EMHEd9EO3IMILX4Xai+swscUjCWZLKR0ZCtS7amVKXo4pqb/AiE92KVoHZj5cidRSG
z/JjQzTzuxKQarotBzJbunS7rH+Gd2NwmuFE/xVVF3rh8JqkbFvZ9TFa4Nm+QoCpAJASIcbO8X8O
cXXw7fimbtaC5I2cL6dOZRYdDPXY/UAjImkGvpZY8eha2E/qSBdxQu4W4uFfx/hSB8F4HX3rD3ct
wnYv0KX3k5/lF1z9EFkSQtPMgvabdkzkatVvX0e1IJMRinzGBZHN0Ft8cTznBmbS9yfUZJhOVJI1
t5b8W3YKd67X+8+hYO5pHoeRTulHoHXMQawYI6AiBuLkQ3bO7WXg0IuuN2eKGOO+P3rDZ0ai2H3C
jQ+LD84xqzHw4JK/XYecq0l9He8GKWsHUdOpTvyvYaBBSkTSRtc54yaiVm7Ob6p+WnWiKr7UzAC9
GAf0CIzyGi39YvdG+PViiOc37GWwyFkqraViQ63olbYGF0Cl8etqd3JoYEB1lGDiQ+JLZ9lp6S6k
plrTp5jOQCk+gOJd1acX4gMkVzzTt7NLdN7XBcLBbaj6WADES5llGHilZSJ9QCCmWpx25pyS4kP/
H5eqxHU10KAfm7HQIYumevwmd4k+Iy11kkZGRZcKvhfoZBLzXCpMRf+8pUSbQ66Nc9EuK5+qve7H
vwN5ViR1REOO06xC2OJNiqMQnoXBGhPcF79+ly6ZD9TkVyP0H5olkWK4B34lZ69WRBXvKbO3+E+0
qQxP2LVzAr/DF39rYRIcFFpoB2xpt38GsvkOFfjBB7sJ2Ul9LirjYEW25VZSF76QhcYh61eXeWkZ
YzMdPgezPPTZ7qnIfaNxtSLaTX8VPytXv/ygYY5CtB9lwqUHImOiGyXZ1osfk9JPUpd3lr/rhOPY
9v4RaLmq3BZHWxDyAlsOUOwicUhJcbU7yFD0rPJgUFd5fFnLC7FDhHr0n+bIOsSUSbnVgXceN+Zh
3aq4flPBw8IxIXoGqOYBjqWDwU356BQ0CRv3Z1reZaQPdgE6MPJ3yoF0QLB6/AL4qlgOC6w2LRkj
y+/CcSD1CPvL5W6HLL+hrsPhnVTCfsISInM5uJK4PszvSDCUTQnt4LZ51WaH/BG+qRCNG7wBx8QJ
yOgJ5vlNfz2bfeGNPKy3glC4XXoZQhtOh7Ic6xbt4n8u+NRFOs6gRf8faxJNX7uPWHPTUiY14p2z
H27bwNjLZVdhVtkUujuSLujNE2walyn8vh5PnE4Ob2v6ygb105nbXLjND8V5NyVBwT1RazgGW93U
B34fLZ0WkTnuSwrAcgJ9O/eG+yV4w2LJyL/XrWDBXlkGddsxH6NyWxcHPeMnt/nXc3rwX1iN26RK
5XKU29yxSdH9y4yD9gMDMzM/WtWQKxI+sa53u8R459MunnSPn9irr8/YQAxHmGCt8pu/omHIpuIm
YP8xirfbb4dTJj44eKyHuhXd8zgYJg3CF8Sfq9Mw3cGTWUMqdkZJ1gv5EF5x09e+2xsJhVZeMKgs
WL7fVTTBLxwzrTCOG3YzflvGbaB+vK+PlhnDgdFIK4VFAm73oSpKoOBIBHOvU9DU8eghc/CbfTOa
3QS/7An3aFUbPtF5YWrG1513pp8cxT2fyLlfB8TdXbC/0Rhi2p0bAjRM0F/qHejh7y+8nXvIpq6U
w+PtC9emAOuTLK9wOXr0kXjPRJqaQzvHx0IV84xXsc8SwerrH7leQ6/XxRR9lrQaWU+FzWemLl7Q
JlNu3i3q7ZVVjM+E3GO8VSVECtiUpK34nH9CDhHDvH64ziQYCj+X7h/uffd+DYgOzb3II2iO6XPC
Qph/jwrMDnjO7Rm7+CKaaQ07hwztydUzfg3XRsDuJUPhMt2MdtlWCC/ljdVJ+0ipH8nvXtC8ZUjj
KWophGi+7DYgmeDuSRKf3lieT0asUkZYDv5skF7+/HrT5CT5dMV9NbaImXsGSn0Pvc5KbWcjf+Ly
WTpWYFK9+OoBRNyk2Lp1nfUPhBBykGaekObdBA/FidD6ImNn5FZfjXLxWBB/RDLgbbeHa/uy7ZbP
5arS3+Ig800Xvu+WYGguYQQP+hDdJO49OhYG2o0GpfnvEk+Y/MlK2NVuCDoA35/pDGhcXeXcnvp9
s2oSy7B6KNBwzGKdtxGuHaaK8oOEqaKwQwKZQJ9ODUbifBau+XLCa16xgij68QE924hb5o5nzN78
T3Fd7dFp5A+98BvPAxuKJpi0GPBEB84MjPss0TKUZ9PfgDwDWfJcdehT0IfJCM9fjnWJO4qoyVSv
Ci0CpPP+RgCQBkboJYAuIXIXeYqYGBYQB68t+fevYc7cyeIBn6g0iobRgVPIHtFAykpLC/xGFOch
hM9/fEZjqnuo4Hz6K9FOzKOw+sIo42cofDXZB6WZubmusicdPrg8zMwh7qyxMPtzZaxog4dZlZXW
IJCpdJwDiBmoo2t8LjBwcUxrURXeN+INCK9ZVJG/+uEHGqBfWAPoRT5KMRPva0bEe1zcPhnftVbj
tBnKR2JZ9N0ByC2Fvx7RR8GQ56zGkgD6HSJfRsYW7B6X8dX1MN17zYAjyd50Gab3bWZfXNnM0Xcz
0ahI+ttdhJBS4vnbV89DNQwP1RrQX7D1AEaRm8glcx3ocqWJjSh6c8YU7KyeNnkSsF7ERN3VrcNZ
pp5Pnsjyos4nLZnATpmW2NRslTfLmzDTiYC2Sb+XGt3L1+I2WdiuM4+ggnWfWOPogpxGz4anS3sQ
YEZ9YRQfuj1hHc17ISlToI/HHrsfqUkXH3G+qAXFTRUgca0owcM5gaIV531J3IBdHUFhVmaSzYfm
rNUs6DvsBRAshR52VTQluGkT7xlkTWsG7BiPpIlRHhcQZJXCkcMDhpCZeUMK9DB/Z4sZ16T7pIB3
wltOQsBIB9WM5kEAQ2spdLG7xGHsnqlzc4aU7kpJVc09qsN74YrYvb6crA7/+jO7MR9KrmJtOaiw
Is4G1n/wtcf9qlsGENTSeh92lI34SDmYHZCKRn40NpdVgwElR1ERUc3bcHW7CPBpqQZ+TSBJBz5c
4aoTgxHnsx/TJ11u2zzQAcdPYY8CvFRdYf6eYoLuTWYFXPE5d7KcurNkUwlGqaotooJ7F9oP8vvM
tXww8dEdkzw3cmvDCrqgSw37q6XzujLetQqhKhucynDJ2Os3p+ZdMAXapfviOUdzSDx6I85o0IAV
QLdXQd+IcLm5voDlDycKMhVp0zbHkrPWAIqaObXVta5dM6V2mIIWG/o1oaAa0dYVsecMhNmHR0Qw
1/iUnNdUpkQ3zIIdFTWmQ+1k9m3xDuTeLja12jQGY4RDbPwfWnRC+Jvb5HX0S3KKV9q140T5MY/Y
4D3FyaLtaxG+Yqvjfyu8nOT4c4rDHxz5slm3SjibHY9t7LeBbR191aIFqbWhNpgQYZIUinjh/vgx
oDnFqNIox+gV34Z00q4WjlplNU4OvrXcmQwAYUmLcYJ67YOY0dXTZrDjHT9WT6LbbD1rWBHGbMNx
Gt4FJ/7OQ7NVwT96XvxXStYk7y7/SgbLtjGO/BHSPsw2smws3zITmSxjMfn+On/90OA1nSgUzOn4
+VteghLWUyAS3pFjtp3fUg+qf1I94E297kMK2SUI56clSBY8amHxnmgs3NlUyKBNLAB6nzkWotNl
tXxUg5EI+AKEThb48HGE+7eq25ZPTRbc/FB/Tn5ylME7UxE7u1rMkaB+Y56yamUIddj+Zh+opGuI
l1Z3czv3VTICkphamjfmH/G4Nury4msqxHXvC80Hkd3a8ccldNrkVTp+nIaaWZWCdbrO6f5nTmRm
5U75awOlMbhci9NSfAQIToFh6vDwNX1hO1Wu5fKkaHe2swtLF7hTlUp++lkfHNoAkXz5jCZ3HGiK
7rcZC+OhivZlCh5lc2uDtNPXnD3a6d5faguUFKOiBzwET6ddpd5kU7yHaYI2m0tFIwPSxFggzU4C
fZDC2ayoWn9fYZ7oey57VBpqCUyoJmF6/ThxDmAKjajZZOloX35NfHSb0BPRG8c6NOu9AiKwOMcu
R4ElBWM7fTXX2o+brWrEBP9yUZembjnjS3yxy/IMpJhcVzO1kORGSBc7DXOcTJwIS5z8AKjitsDL
/prFi4mDcrz0D1fgKokarf9v7L/fBPfMMeXLjY2etvCjc5EJE0WTj6AySFLHEXLxfcbDfxK4LXkc
KtRf0nCckGZXBH0HcnApvsxuDhNUe5UmngEs54PYcBmG42dEQzZrrd+aTCx1M48zOcykc3oWDqVF
YY4/Kn9Z+eJe7ln3yd7LqO2m9CYCVzsIrRCh4leRoEcnNf16gXCl8cmd/Sl1yX7Ltd25AmM/mI7y
AEsFNx9ln4Z3YiJG2gsHKbSd0ChPXJuYthUzs2XayqRQ6tNpTNfkwDKgGuqDPXv2q53THjtbQ382
co/DY2F+DYxq92gUrfHoHENpyewdzTUrQsnLCONfcH9mBrPLg8O6hB9kq58nNydEp8BkM2UiRbmt
HHwbMYyqDe6o6VCXufaaET0OCl6+HaVEMZeNzfYyYQeXpi+Hkb6mb1JKMCAxGUqGKI47FSzGEK8k
ZZNXFzu7WEBOartc/yJ4O6cjWBVXW7Iu4+mplR/wvvPCxsEb4WO5pBRbUAj/kZ1FfnYFpnZKyK8X
1qlMxefwiZh+uOB4B6MeadJW4JKUTFZ8Cm58OaXO2YDvECR6+Rnt1VJ6i1O/TsFsniGzbTYIG+IB
3yXfQuA2YLrCZU2Px2PfL2VDVzU1pWzG0rWU+9mVdo0g30boof6U+7jJ4xZsXPZ+0DeHsjFzChub
Mf+xogeCCPfmWQNBFOA2cTglFKwHSN9OhGPxPK0e9Bei8tLq0iJ3gXUnLqg7HR2OguefkHwhhgUL
eVjSxckcgqmH36yCcCphlqt/ymPCh4ZL0dFmUI1GIokjJYfziDh2N5Ab7Rn+Im0SxHOoeYKz71DB
/N//sHNL7xcqC4yhXCVn2NXnm/+ST0NlEqQ/1zXFMGjw0aAawzS9VB4qCBL692p5GqOO9mSYZb1k
o0Odv98lhTtN01CLOmNRxbY99oGyXYxMSOc9i0TnswV2w0iePmSp3IpZjgEWrQdmUO5Cs8TD+Njj
ebnOrnx1ouNyJF+6XUEclJ/Fpklf9ywySPeFY0ri3YFF0Qv81tgBbxQRlL6M7s72NtOjjY1wcz8M
6IcBoQ4ltctNqit9lbjvn1jYIHUlvmOd4yTT6hvR3wYoLp7cPqkUYU+smk8WllmS7VJxLmAE7Tx5
eZeGudI089nzhI8KD/K0YAGvrdj0lf3AGFOhoo9LnmI/+2yoV0+jU4jtmCF/AB7nCEjfOpBf6CmN
5hEI+wxjucM7oeLkEtYZjD5ajKoO7+F4QL4y+7eNzUumVLnCgdvxq4rkOyXo244eHJQICpMVLpPu
7iyDV1/6diH6QXb3FpUqJ7CVKGCq3Npam4FICGALepY7t/AGfijcfdS54B2yEpgSVwTHlL0lgAn9
u0NpdUMb0npA5qO5pICZtDPz3LbAES2S6oVA90iij+zjHSkiFRmoUR40omEbxeCYePe0hAwKWYYG
qJHYkEyD2Y+53e9Sjf3KFBXJ2MtHuEqcEkTSO7sBk1tSi357y2R6+oEKgUOxFYx1QB9ZIOr4hg3X
YjEG2ducZurh+kW0F8ky13de3FCeFqSajZo78zKtY8TSVtuahhDI18Bk0aSRkvlubMBCM6aQuWdE
GMDw6sqZgiLAdivbDOQmjEjn7gjKZmVESu1fg1zAOsuyPu/A3FtIcRwNe0Vu90Huh/DYWn8CLbhM
396Z90WwKVoKQ4tShcWea7zCiN5rwlokL6NW+U2V3jVYoWLqGkcbVOsaJIFPlHDcnYrsMUMkL5Ob
faiT0Q+rvrM0/li9d2QLSaHgZJNuz3D3nHy4ssMP9qWwtIiVIdsbHrWGDZLRljwoQewOWLzuSN0M
cZ03e0g8glVgSV0pRHLFU/UwQktq6KNK/ZoGiGTZtUWESq2oVLrRYLxbDg7NNYr4jjhKCLm4nFI2
uiw9LoqmPXuPSefAa5WV0v5p0EXlK41SmHx5B52Bvi546L3Ng/cM+x45jhZtqXusJLNfy4sbsz1K
F1kj1euJfU5gnMscAXL7SyHZWMDvYUDgg002++U7oOsNOXu7kYhkJFv1oXUZBkYdNeqs5rtwUVOD
HJfj3JYQeT/5ppevb510+55JR2LMxIx1Zm8/IecMKNV2Z93b+/u8vYIqGmdXICpu2BMVIgf4Ed0c
ER6jWdzEJjKV8pKfgsfHmwhkTHRrv9ipwlOKStVz3CPV8zBJHWY9u/LL99e9hPg7Yw7f3RH8vBl5
xAxNvagDCbZ17Tqh94AviqSDogQIt6NN08vObuUrpgAt/4LkAWQ6bB+PdVHEKfCzeY6ByUCnAFLw
hqG40RDGJNiKYrpH3m47pKY5SwFovmFg8ePdUwEfBPIt9RcDKgbqJay72WakPKHJN9TTPA5VE65F
crMfuB+vvCigO32JodF+w+Hx+2bHuC6QpQrTh8yoKsVyjyjNbxGhECEZ6wU09WbbIfA2DoqirpYt
S3yDZDG8ybm8Eo6krMKlAac8Yy+SFma1ZBvvwfSb5LN0JCR6JalfL2Ygju0l6YB0QQuLzvxdy+dw
lWrL4SgOYu2zkwJKWJgZsJ9ndcRmsYa5j5Xy2Y6E9zVKDoZpEBA7CmX9Uv9xGdCqccMDCftOeOgY
91rTXQv1FLBuvE198neDLVTqBTNqa+oGkl5kzPpMcWjylrq9JcW68m5sHmXsHAWneqEj4hzRcE2f
gWNTL/iH9JKmJEqp9RPpSfnRaVShn4/U+QMRu3b35AfDrjinU/2vO8REUuwUsJv8JHe7XVhSvKF/
9Ce2FzCL9C+/STf4mEFefmTREH/cPSeYUN8HG0DuxObpfPJ141ZOFo0sfzX5TlWJCEfl9bPUMORw
JRBsCehrJa2jqBg57OLOXg9NxLitOZT06J6jFQwOXvWcBcel11zdPAl65oOg8Y6cI72oT2sEW29U
Xa+J5Rx6jU9a0lD6eNPBcYsuFTuhSCUaQbQ4UgaGTStG9KySUtCa1jf318bCA5iRdVPL30nowIwe
cirukDbgnJNI8ni9/w+LCbXEQmYphPd1sEQRdFvnXGsO0YC3UuQhIDb4RSa2vsvCYo7wSUw6fcTj
cpS2OtpfE2jYl5vCMLZr6dnrCbWDOjrGvVkEN3qh/lk9sZWj84Qb7lTG8x5th3i/Np7m4VpSoyN/
51LSFzoiMrWeBwO96/ziHy+bYfJZU42mEmxnsvadhLOapBklsebc5ztqZ1hy7mCY3zj1OiB+NRV8
cxY634icmkvT3vnVFu4FVYHZ9S0hjPgdflqk56efaquSrlNEohQigBUKIUoULIN9tYADHQZFY7Wd
le071NvGjiiup1Wji264BtGO2gy+GA8Fu2TLLFJuHf75XcAzMZjlWg3PtntRVLfJjsjkHcV/ofz5
y0T602nnpSmGTexm0KuFgX3mhE65dvIOexS4G26TOPA/3xj/C5hlEDAKfNBGua9XXhjy4F7aR/7l
MbkyZuf2ZKMb8BoUpAWO3IbeMwNS1s+Rwz1cXetyqsE8GpBUySU5JsDRclNGZ2bHoBqRrx4rTiLB
FQZCoyBcYvCuaM/IIqPF9j5I8umu0L7rM0PB2CPXHVukIlDqhNuJXltOcWSGiGXii/wZMXmr2e4F
yyQaTeLUlcuxblHypWQN2LI/n0WIjGwtpJC4acljpM9OzL8MfVFvOMPsVlRIXh99JV3EyuZOiR7M
ChEJip2VSCzOXNQGjBaUVGhov5YOpElJIDqXi2DLj06QNbWHeYi/4X28GQXt0f4n8LgJYlDjsjow
Gt+qgmM7yKFkeUs5Wqgm4huh5KcWi4TOjN6ihgza4MS703JOIkad8N128ORfdxuXL8z/eUqoK773
K7SaABALqcziHgYx9rJVGoG4grTqmsuSem5687EBAMNQvdW8DcuT2Iewz5imsPZvPJIcnj5q4vsS
zQrNVsW52t0WwoZw9h10xBcZNIV4Mfu8lIQhYx/F9dQr6J4i3syE791Xq+8NrZm2VDhDgJUpR/Ub
7cpSYBeZB6+FJcexSIdOuSMwAfLbLO/yDFmjDHMZ/clA/htG/Dup1L0XaUCHOxm2fb8c7W9py8Mg
gflyNWSG7fhsiEEu/hdcSnWT8JTqPtmdoyIlFxIj/ciKxjkRP4v7C2iSmjeH34CxmWxMVk4diI2j
MwFqNLV9wyQasl59oo1jEuVJMgFONHpKYheZSoxhZyOMU97C38j2WTJnpuqt/bXXjqiqXEvsJfWz
CwegeXVvFpysrQLgLluiUzgTWm5z4dIeTRWMDfLwV84TAe6FB7n/H311bf5RXeRXBNdEuvnDYL4/
DHYgVeSXY1I8lOwVJzT2rlRFb219ot42eC/WiI6gteCObS+uYxVeklVgbL/u8GhRQtx5EWU+4pYe
6H3y36tZHFB34TX11/t0yRnNTYS+5foKfN5O2u0AKZHxgIujN7EfPeEIPLWt6EP2p0h6py1VvfIU
J7jOnG0ePG67dRPiZTYYNOW875fr26e67JIJjCMznLAZBW1XhX5SZjNtkGLrPatv47xXsow12ltG
UwJnjSJb/v2NXbjVwsISiOMDkKnjriFhGew6+5GTLtySbPpdN9TBOVlqKDlrVQJAKBLqaG7DnYcD
hY1dqljoO6PtRgUWIgZ+UQzyLNSUB27fXnMXaGisWs8cTVIC4pP/slApkAeMchM/Qd6T7RRjgBn3
HV57mcc3oKpOrfsNjgBqYy/XOqxvIeCTYEsmrX+FNCDnwGLLQhrRxV8yDo5P2zvUjuzNrbNQByAN
yxTNzvt8LWJ0IxBDvzlSI8CUC9M5TEpbvHgGASdws0xPzqQ5aSZpmy4PDGy+i3ZFBh24aEQ6XJtP
wZIaxgGrbtJYX3kPtk0pRouKdiKmc6uMoD95XrZylaV+SnlGG+314SYQm+PBYxi4JjV25m4CMu3z
g+k2GceBZAX/W4m/u6misw02y54W69oY63Qd3skkBBSGSIdo/761jMZNoW1W+6bcUizNUyw/Jy2b
OJg3waEVZUJu/IsIP7QDWNmKO/FqaZooAALZ3RWsnnofpenHooWe1781+r0nRwxm0hKw/dUAcwfE
HhZBdg4hgUv5rN636Cqww1ZVHvQpW8Mu66jNqmzD2qZpnpuiJwJxpAkwAt6Gx+o12vw897+v+bQ3
4teMt4rmc1EfnOYxbXMwi756Ma6h6vuayvErXVVwOWIwCwhi0L+uv/Vy2Ct5CZ9QaHEqioeICI5+
eEhlBlHHQz3Jymgb74P3mzoeYSxrF6UxNVzxiENNjgLrcDSxczHJkFpOLGA76NqHDU0cy9c9wHvX
1eH/aCe2CdVTr7GBLQMw3Br/diKMT2SvKswpadN9IBQQRGIIUpGrThY7eSXwdUUGonNfaFwiMH+6
soEpmtNPPVPpVMDGgCC6wmII+Mc3j4HYEX6yoyLMT7pnlcjhqmrbi8Qu6L0PlzinW+emUpR2uqVc
QecNlXQ0at+3YsPoGwnHMsoW2yuuBu2Zvyf5+/TbJeaI2fPML7PBDRC71CyvS3R+K8RIMtPuT4/N
E/pfj5ldQZQBmv5I/Kp1JSQRBBEYgp/v8LFaGqxHjVHiALuaJjqyZagBSQXDECRHbmWWX/9+y7B3
LOjX99RlabcCdWrM9+ET860O10pKrQV55KFsIo8jKetQsrMi9FnUo423UR6SS5fiPxaRlVxDOYR3
keZ7IKvhcxAbTk59jYLuDRr74rtjtwYg8G1ViurAW0lvyTEf+pHMZgLjx/C2cxykktB50bWCIjlB
cY+ol/9GwkAM8juelJKQDV/ZarGCDPrz0AANOBqIvYPSloU3rlZFGOmB446X+f4c5molQK92rRCi
xdEPLxbIsKhuq/4tZAGxCEy+EmUpzuO5OTzOl3BV8ddlLnwVCBGAoLGMfT9gC0onTBrLFgD/3xFz
zAiuaLnIoc3RqXtkzJiKi0ags58WnBylHST9rf4u5Jzvf7O2is7SANrP5CtF05etUu10dYq50foP
dSQ+ftQZ9pRWnvQ/USyhcJonTs9fKsC7y2UDXDnBfSNCsKnkC7zqN/ou12pjWD/PQAHMN0Kjny0W
MvUmol+MXe0D5A7qYLn6MTwMyQYz0Mm5UFnlIpZtCHEXPxx7E9u15dVrifW2egZbirei8TsBdG1T
q9ohifNEHDoMINb/F656X/cxTaX8o9ynCv9U2iGCPXXEqNhUmtw/kaJbT4M+iXVt01gu93cMhniO
Pu1ypC3z0jv1ZZGbZ62Eb/c8LGLjuViREhRW9qxGxx22Rlx8ceWLth60sp62VF1Db7S/WT+OXowT
uSzt6ZVQp5ni3Nq+jqy2xce1BKzdnP4rbTeHdBm2sXnUodsDhUoV4k24FG0N41CmiabHue6zheg/
pyV6yyiOw+OMAkCsaig2M0i7956PZ4Ot+hU14kiplpfseflEz2E4MLiv149GTP16cdYN3DGWZOvp
jh8LWySR/Vboi/rLvAg91IdKiOGPqKKUzFk9K0v53GbvJIXh0UquXAfL8TG1lrgsHJqBrmU3yuLN
LRieNjCcrq9MPTKnGr1v/Q8pJ654iIk6wtHxnYTrXLWtRhk+ECRmGN2yqRjpuRjbd1mVXpvvC5FB
9nPparyURM0r/pMw9gn7syYGUA1q6cK8N9eLplJsjd3+cHQ1Xotv3eMde2JF/cvomRsMyHbYEDGu
bhmP2YZz7ChuplIuSZwv1wUn+m9FJMLDPiKirjHWPwGoISXnSBmAc4S7I50ntC69efxl498mXdeO
z86oklWVjDZFwmC70jt+3hU94+MTzS38Npj2XA1Al7qXEB26H8kQy+6Yq/BOSd6KIeDlstSvJ9Ln
IjiZzD0Rz/Nc+z5vSFRsWrkxYmpuOJ3HG14/P0linA2rUYussJYkBhxvfgGEeeySMQzmSxOxqPvU
0O4960eiIqsBcaYKKRQRWhQyaUNbgJr2AHmLyHXIrnUaKx5yZ94igcxqKu882FkRZIHyeB0Dasvw
Mnracgc+KEKuoeQuZM6V0r/G5kkiFct0wIDVhVzY2rrV486RthBMVRvKdMdJvbXb9iKoHDaCUW3H
Su5VLfZJXu1jFPsbTp3mqF+3mW3OlTL0YtqABLcdHFkeIrM8TixQXBOtwwDASPWJPwS0Is3vA0i2
9rhP+NvFBly1pWAfa0NkWQTEDsJU3RaEX7jV0VQIHbQtw7PbkXAF9FrYLoWul854SpghOEZ+XKw7
7kn9UYGs4y7+SWQr7uwToVcMQnNCTgjYjr4pHbdfrbisdDf7uORiOIZO1fIGdsx/Wnuzw6nuU1Fd
s6hOCsCmYHSr198hJS5hlDdFz7e1zhXjpRjWcR6MkijEbvOHWLNEV6CyEr8RmZDfs0bzVsCeZN09
YjBPtKnfC02IIjKR9qnNOVeBKAtJKwQVBHG4Q4gAREhF6ISdzItwihdPyEyvNd176puVIGJ4aZjl
10m7e7MaoEto0OakPKiBvbAT7uV1SZ/T8DnsaB4IPbIiovZmJ4cjPd4iyVEZqEKlPn1MeDeer6cO
d5Hu7V0U+gMVH8UEc8IvCAwxoVdAQgr8Zt5ncalSb39ZZ2N4ERgeQzZ6msn/yBp82lLfOnHIEhDA
9MfjXJbeTAXMjgNAT9b53uSS9154Z50usOp4ev4sh5go8+SKSI31SSQNTHcNyiU3iDEtgDAsbemH
R1R/0C28whw3qfR8yDnSF4GBpmSGdQuP8/4nme/ux2zcBVoRv6Ok4xM/+tBViL1jsMK2fuOHWWYb
WY8/8fzW3jzJUCWBjaGtWW/T9ZVesp1uyxxns5n50BLsaPMinQItqmU4XvuTcZekLStqdefafFTr
g4an14iFFZR6jJXDYAkGezlzfpRtWOn2hwGNzaU0h5ki6tm0TlBZV+y6taLqD+feOdJEU1Hkn1vV
eAFpvJTh5xrfXgW8yrY7PV9VE65u1bZnjWZiWDE5sa8V7GFKy86+WF4AaLA2cr6aL9ydzrIf+pqu
LqGpW8sxsZRgvJR3RZyjT/H2eEITX8sdG/c+Pe/2FZEX526gPv3sCky3xjLS2ao7iBIVQJIS/bhU
H0uBIDtBRhawwhBZQZ833M+dKzPup2puhDD6hLkmfKA4F0tz+doX63QeOZ9IgrGnLvOG7zwskhDV
AEysdz3Jt5Xu7O0cuCL85xynqQCU3QcPAFfadCXk6n90y61Sa+1uyr9IYptXJAIYHs7qTkBA5zc3
x3msUygDoJl/gANhrqRoObbnCfftVDtcH8idfu8q7thLluzSqKd+6lL/zDyjSPgmkFT1IZQqfXMk
QGBpsCjfhOisJ5AUgZy77Xja8ChkES0JxTASORGo5awR3M+T+bpA4JFj1qgESeaGJiSH9Mz2rUNc
JYXgrlPdylVdY1iSd9ihXAsOfPZq5xqChhdDkJYiuxuHjMPaXl3dQuTUK5H0+wsL4KNXBcCr72nO
jN+mrXVoy4GMQLE8ord0tg/spI5n9NNFMWvoAAtX519d7dS2lBwvgeWuDVR4r1OLcXYCqf61Gcrb
NNOdWH/IgyZMtczQ80iZziPwHF/T9R7bcBY18Ssc/cGl0QGC1s0KMGdOTbOUIwu6L+sW/ldBQRS7
Rt4mjdUGcxmsTBd/4xTfbDFqHgAl27sjESshHLbje54vB4D4Hx8EsO/tCxiy2314QS8RBspU8IAU
oveQvwN192Q9JXJNhPevWL6QumG2pBu4oUWiKfPwNvy49bd2ef0X7uYIlLEqsh2F6zztqsKblgzH
4TdNSZvjrme8PKAggyg2F6B+j1uI+iyVzw3yl1R1A7bWg+Nih8N0UG++HYkl0cxnOhnIwIfGrUb2
TqLiV3JTJ1LeFOkstmnw9pYxLdUO+Zls+/z0cK2HNQRCpq+0h6WthhBDUN7Hrp5oiXg9c9tEoBuV
QTT0uhGguEsiSt513KCXFZLdhlL1zcEMNH8gTJHDV8ZnZMCO0Xcju7Qr9O6n0l6O5mwcUD2EbdhG
YR7UWPdKPzf3D9hGcLKjdSWr0JGu5O8ab46PwiyKbBkodBmcD1G7Mv3mN93ncf0EDSCVSRw51reQ
ZS0kT+tMThy7xPvFu6jGvDJStOtEQEFeRh8920gUsQscW1tGTNHyVlYTWPJb8dAkXMCLijO/sULt
xtLwysNsiTL9GFX9WVoCewHQHef8psHJ7VT8mNHFKokQdi0hQYIxhiFFpjDiuZDO0R08JjHixHfE
6lzTuWQPSYVlZqAFHZu22w2efj1WtBGId8RO67Qtb4A+klhORLPqMPtucmM9C2HyOVLxc0jcI+FC
zRKS9SrOXrcg75xBptDabk+HctcHIZqBcAkrJPmSM1fOZluz4KKCZcvF+MezMVk8jOc4PyA7R4IP
BFgjAE37RgjR5+msxg48K6xOA0k6AlwyZOZoZtjYmd0VnvHv+PQhrBe2essVgCRukCftz2j+DjYg
TSauCqZidWl61jwGJrGexHDO1Grrg47wduV2wiOH1q+rBi1yedc/yV/aZhoINtSHwTi9IEbt/f9x
0Qb2jagOO0fUx/VgtwncFOpkXB3oIMEmkqk1S9wxCeG0dSIyuQjiaCq+8QawqjhU4Y6NAXiftW4O
6Liyvv9wEq2mAr107AIqikkUKJU3yuGE4msCmsq0h5f7VfYcHl2g02oIJcWW1u7gcz0N8SgvQGh/
8rv2GQrIrAX8u8HSeXAti5FD8K/3ZoJBieEr2WnLdg73IyKlwnb1WxhuKO5O3p5RV/ncAFmzE5lr
nnJAYyuUiEyKWHiFNCR1fem+MvxShUbgeMoh4OkwrptZ+RLgURcCIFHwdxCxg80AHCpdpr6yJ4z3
Ch7JKgPFFQlUZ2Ynl5/5r5GpjTRgZMb6KOlRXRZ8W6r3qQ/VXSQXdFrzTiuYlqD9EDn2fMvmGl1+
6IzjF/ec3ZaBTJGqmdih3NphNJKj36bv3xMqTctn+TwXU6Tbqm9xr/f5aC13Ci7E1U6zIGwq/3eu
0zgkxuMKBwMIJuuSpLa0nu5tgxkSGcW7stpV722Nz8b0LBElWbvxJuqH0n+++2bl485MyCK6ofBj
3wKZt3EG2C/79Su4sqRdiXaiUXH1NTS+9o1r8chMXgLPVURxG2qi9a0j8OVdq59HdzGvcuh1E/OQ
baxKbSSd0y35FtlCjHV5My1beseJIe6/o7nl+WkoXq47bTmUKcAd92s9DrcvEpDYRftPuBcHwaTV
bfMY6AjHleqGtHoDOKJQLRF8UDudtaOGvpr2mF81G/gYX+qJJwkglUd17nN0uNexksvFXLj5CXzF
1iELfVNfs2sc1ZDexKXv/LGR5iU8AUYY629xvkzeccMd7JzTUqGvw2qKApXbX6bz9C2DvrKklJR7
K1hv9VTyHcCEra6jfH37o8zK1XZchMwTLDAY5o7+6ign2Dme0NbHFVNu4CFK7KFc14hV/VQZtMh/
LPf8xxldQkyiGpEKu9+xrg/xUXWpD4er0hRA5BP0dyDGaBosRjwBysO19MxshCROs0T9e4OJXhPD
8Z0T0mnQo7iLvsX6E8XCF1uFNjp40Bpr4Pa9zy7FfMr44VQnEGFYXHhLpUiuXAqpeHhep4Elb6yW
9Si/BtcvAp3agqAKQJi2irgMxl7vmrV0MW/eDV7wlHeUjfUqHROM3UU4DKcW3v8179huWGnszvLr
1s8z8phrMD38BXyxsgJeApp8p2iXHWBTeBm+/b+UvzfwftDVeA7fFnZ5lR3IKy2egXbLEjVOi0Un
8jlU1JsbG9p5OAUuG5/PYqHn9e8Cu3AYlqJOnWGhiEv4Ea7z0e9Dpe51ZX3K+5qBw0qmqWTh+uSY
Imx5WOSH5zJLiiLbm3pdZ2kHp4psQh5+TyEK/NKLLnFZEiUn9nn4oFW7BSU6T2BIKM18rcqRUgO8
16U01028F5xJhpIhjNBDPJBX+pUcEGTU1mTwLWOboZkZXHqPqVIcBlScRToDQoub0BnsduAsTlSY
h/UDD8iYOIM7IINLJBb6iGWlX/zxDef9IQ4CzkwD8SPYViTlUE1qeqJ+VE5av++EwTSMX9p2JB0V
HCUjWZHV+etHpPhG1F3k32jLjjQbxtAWybRXnNguLzYkImwCoav2UDkSJvIOsooAQsXFAXiFuTVr
9mS3U9OqEZJuEywQJXyMuWPFtPyJ+JEgdYuXmRAaNrM+Dbmjws2/HBnI+1GGe03uN9EotU9kXxO5
FJ1CGvM2JMZw2SLq0iJL9amhLboPwX7xW5DimB/e8/Ym9IpvkHOifXCARPGk+CvWlOqMNJDQxZtS
pByRCYYSGndWSn4Z657KdA+/1V1u0Fi8+58X7NphNy/7ju0ihrwhTmcwlQuagNosQavPBNhv1oET
+CuD4DhGWQXZ2jU9IjIdeKjxtDWPhTOs1T4NVuaAxa7iOrRzEJbh5wbY1dLXE3PmUuw3vOsmADGy
w4PZ3f85LOjXXGp3g9ozTQRpri5ch43q1mZjihcO7xSNJ7fjY/3ZLfADGT2Rt0Y7NVvyNaG8kvmN
JM13qzgin2TYi03Rlghb/Krpi3d3HuxoCnJYtqD6sugFfGtTCJbDkUsyJoHsITixNcQ/raSMa4up
Vikw/8lBngY36PxQuRXdFJ6v8jT9VbfdFHKDRhL6Y1MoH/A35O53jLKG4O0uFwgvyTxgx5pENpu5
mmLvnXL8fVbyOaojugdlMCdS9clZlJWPYSQbDEZoDEmEHmJPycuUVobBTRNifw5BnjjzG9CylUS4
JAOqKEKjwqPLjtcJcQ4xoL2SnhqHusWh6E1F3DkLl4kGzyipWgP4L7Qsu8fmGg5fU/XWdpJkTSET
C/7ds68Ns8r58d9j0whzi7qAJLUGCBjaAPEyzuP8y6g/8KNNj8bgoY0da0uK3BdDG/u3pXYa/yNj
Dv3D0yKkERx7PVwzUcVie3nUKoYBOhuNEyOmEdqDONuSzbBAFawext1iaQ4ZSWfXXDZhB/npqaBX
ld+ubHoufhMf5DJILK9ffxOvw+hpv510Up9izC6cFPEj9LWJIAixa3dDKSY9+JZoGapqtkaVonbP
u2qubwbw7kLNvbzZUkNNlls6U40E80KOsvyha/GCRlCkn++UXTwzqpdFac+iJAm+t7vHMWR28mvV
biDkyf6Xg51bMGEjFPXLnqKgV49VK2uprl0j7g6bxn4eTKjHO7GZglwO6pU3HJzXs4vM9EMi7+Rz
cPmyP3jouiuNMnd8mLl9Bd+GFaAA3ep1IHpqhnDX0dTgTFp6S66w4SWe9T/HzVcifrQJLl7bNOc4
xudf0q9S0lU7n8J2lkDFU4NOpgk4SRDT3hcrCpxcF+nNqdDYu8p9tIUb34Fi/TujeDZGEY9DZ0Jd
oFwHWt5M4PDnb4lkKajnBY9vGabfVkhCsycbMpYcGXK9pI1Jo/9ROEC9EP84mAJQYkPscpzXcG2/
0Do3pOCaQmy54CLeBT+VQuELLwJ1zeX5vxjdYalMqv4N4dC3jUg1E/VIVNlU06FlitHpJEIhyk73
Ormw6ThRN5EXunwLHOUAgyoS4hMTFkQNMTTyv9IlziElLrW2je1MZH9B/u0xKHEgi56lY1tKqvhi
lBdDGfEBIsTWoectBrm8Ai7SslhZuWYh5VTPoESmnoDLor8SqNA5HqO+39kpzPZAYKdDUT3Q3wly
FTnupD2daZKazqW4/5zdkv8gVuUYHq/QWxx796TwMMLdF0nB6JSYyxDM05mxssEeGwxTb7CoyB0Z
Xf/9lnJVYNlRvCjyWDPMhwn3JvkWF+DkQ6kLlcAJ7PnBixNGBBpPHWr02RHyATF1AU6r5TzI7YXr
bOKucnJcE8EduKH/tZp7RjA1H72DWOq+ljuOHJWccJj/yl6n7adS7C3Sb1HRJn+ELWQ2hlbNLCJ5
vOhSyDfDG1uxY6rMnnlpBrOucH1EKOhNS4GXcjncwrQyoexzIjcCbolUZ/9w3n3azBVDdKNj6Gw2
wl8JfDXToxJsZ/N1SeneZbv37wtlVNDbSJyvNGQJ20MweAWZtsRV/64q+fLQp72mxx2IU4gFJclc
FDbTQxvfgF+FRsUmm/lBRcxODIy9XkcjgYf1kPaWJmBCV4P3f/fwfrSvVrtRMV8uhUoBjZNGuOgV
75ftPqUXemB2F/idj0juooVI7OzglmtF5mQTHN8Fs6w+v01OH2sAwkMZwSFGrWbJ7w/R2pH4Yc8z
exGqH7ahhzYSjXwTEVnYx6TvkgYKCdJHhRApOnMaQ4ptkkZksrMsOh1mYLrVxK/FVS6Jsg9cEaYj
YFl0w1sSZlDDc0VN2MNJgcIeMO3enJx7T08PD1ysr9CI2axq6y/+o3KqlnQ8xv/7OHkIjvI8336H
5WI8EJj24dPxpWr/4z5yT+siPCZnVBsyVlngzf25O8+LZdgTKsZJHc27O/1hpIRByPo47xLV2he+
+PLIMptBby0lWLczAHYs8Y/3QNElRNo67X4bCLMbRXN5JvZBekO2M/PCi6fgAhmj/m/sP5KPlGQK
FWh97fitKQvgww3DkJWtVfEp3v2bhxEzSJn4cxnK5LiGnY7rDNf+yXH5PIypgzbvMVoMnrmg8gpg
5LkUBS3hZAFlxXwPlKCZJsxVurjWiJO9DxKlck7d0dWeZaxluPq76N7jng9ws00sTrAIHoUQkdPO
E3p0tvDkROaCzFU7TU0ZkuZ3Rgd6C/W3bHYiNjm0aBowNNoxNYBGHK8iE5jhZuscS6kBPWCn9BgO
96hVHHskmemLOQQAxAuucRQIRm6RpfalOE6b/3SgL4/P5N3zbgpqdcj/eVVtRwlg2BBts5d1DYMu
c7O1ZN/76hvjIIp+yYbys30PtKJRMTPhoau3tyzSCQ02TpMxCw0yv70fMgK6Spgnsvr7D0xMyKPq
QII+n7e470nA8tiEuPfbVOg=
`pragma protect end_protected

