`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
cWZqnfVmlFHGMsztW0Hoc7/jv13IKVWoMcCSyfX2Rb+moyruhqM32yrGdJKnKnm9lNCt2OZi/EvM
w6/MvIMCSsq+XyXP+buV9U1QAbAU7jjnjfuJuLWILgs1zbK63qXQXlNeHfS+RUdNViX9JDB9C1Qd
htLD6t5NN+8Xa+TbYLkY9Cn9o+qcsVBXYO3puD9kMC58MkoIapzvSOIR9+Z44/F5fEKAgvGWDEc+
Oaq0alTsvzKEPnANDZCJOMYQehXcjX3Vjp9ISrnkuN0iJPcDLSoZFwgc1QJ7yrWTNb7Mnbw0Lv2R
ypGYDGAQNjwuHZ62bXgDJCJGa0oPAKO/H8/Luw==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
D4bRrbWQHQV5EWZhL1/IsLtn2FIE+0yhJJrQU5GrEGAzfNuqJXPRozVlVUGDCqIJoPob62eaUQA1
wRIiU3QYxFLv40pu0HsfPWsBD4J6ZLjt/WiKS35eolRtoA1jMt9Jrpr7wYMjbmMOGKi6E8OAzthv
8FWY6CAohieZ92ffr2lqpgnIMOVK6rIwVD2hUS4kOsaZVdrjxz7p5uNJ8GrdclF8oxbLhE/5vVQ+
kJ6lxsVpouLBiP18MxDfisYhKyZY4nj+wGbWEx+nq3UzdUXSsnVeAGXgoEyUcb65dXXb6ZE5QTKO
EH3dC1NHazRiqzVmml7AO/1v6LuVO0XTCEazCAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
N55mId9gWjY8o/vpVggvL50LnvLYvFlFBx172tnnLcguXaKvKNWnMeAzQg/JJLRvuyuBzBt5n7Sg
no/P9jbiLQ==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gj7dH/+0bZhuG1q20KVmjuFQolZ2wLgP7GCRHO0GPec3rfk2FfdatX+sW1gWiihIVpxkmzNQa5Cy
7syA21ZVB6xBa0yaCMc8znO9tScSYyy6z3V5JeyoYRLprPIiulyQSdLK80ce4BvJYnJGjDkI1mgk
T6DoyNGQmrjGSKltsy2ekXMsBG33VQV2aPGke0KFYBRUzRZX/Xf8C2CSJjY/JgW3bMpANot5rKJK
ucpiwetvOsocJnN1MgrwAwAE9qdDoqGZcxtk1cS7qShjiJmoW5+cQUOPWMStXBUSHzQBJzFsRJUe
RjOvC0vfX3kOx/kk79tbdMle893tL2zCs6gDBg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Uo/rtmSYdAd29BuGTO2XaLGG42+mEc0YWuhhM4AUzHUDXnSMog9LIyHCIYk1IXvfyb/YnrVz2LRb
A5p7Vd9IckEpr6gEsQDZkKX/2GX5OJ+mu7yjJ8w7dPWMzK4svm93hKanv+WMX42YDFpnE1GTf8St
W3mU4dSppYuStWGuxb8I7SRw+ZBzH4vwXDceJ0Sshqt5hE0xPUOshwlDLOeLGqgXtI5CtZ7zyH2h
7iBRxO65jA1wlQrZtigONYUy6CIL0OvMZz8I3zGgUYWIkFTuaD/YRXgDp1mBPYIu0vNENpc+MhPc
ADxy/nd6tGnWnpywRDfa6/bc66wuLHgxAEpesQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
A0oc+oR2dyUg/GWv74V/0deM6IbPOMLt16lwRAzCTK3iGV79coLBnDop17zi6gwrojtsITTqFbZp
+2dzkcaqT9L429taeNQa+WOaqbOc/faj8Rgi7KJO86NRGoDpsS77toOsFesNbDxPFXIm67cL03PL
NVLlKSUfDVOXvwL7K0c=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NIpPZ0kzT3P6KNE/hcoIjuKF+zDeW4wLolhaboev+rwseh3cmaifBzTtgC1rkCvFu3UrBejDAVR5
zophCPtB1oHEO+hyMBz9Y6hE1NY4PC1RPYK1TlHryZjDbMnwOegpZg+zfvSrVVJypLG+7miHW5zg
JURD7lG+ZI70AcWNYvjKTILIkO4RyvHoSG3Jg+wUWTKFeX/4MZFqBZR4p2hvErHvswjbihYNNKF6
1hlC3UnInba96hYmCV8jrEG2Dmg/k7tKeSiCkTN4mBytZcwdcsptwE75xv4Sv5r73W89PMOaHPZE
fUD48VERuEk5yLPUx/ah/gwT8XKk717rRh/H9Q==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
uWnwhALj+ZGs3V5cyWMjW8SvO3O+CdtuRXNTWgLp67rRVk2LyHGG/K8LEMnRYdyul4C/8CQk8zF0
fXKJgPrPHZxKps54CvPCFwE3lP2zrxX0d2NH+6b0AMgdNwT9WaiBd9hqj7ul95K1+jH+WYvRTAUw
4x8Mh4T9CQBTDbp+78ugQPWVOzZoB5wh7AQb2wJI3FXA7qJ0FEXym90T8oAvrqgFKFFwerWwo4Wq
pBQdG8HmaIljF3+RxhEXDftp65YQsCf1Y5uLdMYfQlxjZJnCa/5RoPrSgbh5evBuScF4BizsVbjT
rp536/tsEUCJEHuDVT6IvuAfYyTSrt3qouds0w==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
sUTGzeyJetISPOc3dB7p3IfoH/D3+sH9QaPxVaAK98c625Zv2iaOyZOf5qT/6Hn02Rucw5JvJu/H
mARiVrJwXa85aEM4ALAcxFCSXNbC+TqRdaFcU8zcTtVTApFcFZZI4X9ApqD1XzJRCtlkBso45+c7
hCQSCjaqH+LPpovQMJY=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
oRks7kPaFGgS7Svxysu6EGesX8erOBpeUcKUq3QVUj+FOBWmtIoCDQbwzDsGjX737myvdVbIXyqF
apOnT9gqtYCZAIMhIL7kkRPMUXUkurs26y5pylxE8ocZOw4wQ0wtltQOuAM4EGDKQJ1JUrJhKtGP
F1k8Pqgxy84Swx03lxdgUfVVsU52Qt8NtYJZFu2yYMFSTpXClFqTEC3UnaIJ3rZc4XV1qFZkWnBR
JHtaXych0D7cqbuw+QsbGZFyh2/iE+UEPxy2u3H1Ua6f+HWeYGpq5d66w4ls+O4PYAA83WsuLXcB
9A5ZLfuRHLza2W0GEYTYzsOFBHuWg46scVHJpw==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17696)
`pragma protect data_block
9rXtrbVovnubpDZc+edvHFbJ7eSiTYfT/3a7kqJqoM2mp4fGpWtevUyr3a1QFFmaLEsIlgztupm2
z/j+52qVYEt06ih8z85jbrrYu6e7qY5YPqx5GvjWC6Ci5IAtoM+9aOHygLyYCpiRNl/B37asePY5
StpnjDn5yIuhm88T4amTcDxxooYsvXs74EknLo2kUBauUxMic6EFvYdYsCn+DX2EvtWjCK7hekh6
Q/VJ1HmTl0D/WyU6GJ/SH9rg2k/kdKIAgvok7MPerUxXC7KBnhoL33OD1TOZx3qoxZpQ90Ub1/CX
3MNEBEpuM4XyEF43XbjvoFTaKAJxSnJMFxJ/CNKv8kIDsJmbBgfJk8P2tMIu71tKOGTCS7YIcltG
6eG7cNzSbR+HRdveuPXgAyji/Ozvf4Glqkb4zrFVbuHbZGE9yGD/uxmOTIP98POV+soh61xzUYOB
LLK1WfCE8h6c2DGyFq3DreEofpnD9x9hmqcS/gLjMT9Wec5ZtZ5UoGlqyfTQHZwhZmLLeFgHsrr8
O7MITMFjjRyMoWOb0dWfep+/pBge2uz+I4MgsEzBC8040GMp4MakVNApPOrNQS476/uqt449G/ND
tyjYivbTLdNWHa8rTM6u0Bbayb6qH1zRqAKHvfFYI047bKUUXGCLKSWjy1NVB2inOut83hiB6M7y
V+zRT809ZgpV3/iR9lPNztcDwqfzZaPBSHdkPyKgMmUv+UQdHM+7EZCDNW8BCLvXZKrYLnF281gX
bauaHNNO1eKInSFY0SyqWn8GltuYrRaklv3N+B9RAqEmnJiE9SSGXRhBJw/zyr8bPbcb2FTgfwSt
xdo+A0LqsKYBctoB6shEAiB4lXZyRN/eC15nqSeiuJ0Xj6CCfU6g0XhSzahU5hFHIwCdibMRyRAv
uKV4P2hMJsVaXraEjTXzPV9Z4qGRhL1zPgiwNX5fuKiQbkIb+VQ35b2a0jS9/Jh1X+J/01WVNBBA
F0yoXqvcQk6qb3IPawZWJcqgoySTryZNxoma112FhcUcJNpGbboVHeBa0SZudK0LzIzPxXqIhHUG
m2wbBVDf/cbP8Noy2Z/FrSfZiA2wyTqkyvAdu2x2NDRjbZuzbP1QEH0J61ZCyjLjdZ7dj63zVXp+
w2jx4dh7DR0WePNPpNkYQiy3o1PvBaNi8bIH1FrRC5XgYKOJXhbbrq3xTqzH0g9SjuWTL1MPNqB3
wxS9/w9R9mmexUJchROrpdkrKSMviD3ZDUqpnvzgXUMFXP6gZqHvaceOpsE29zJ9kUhlQIa3dLH2
0nNzeQLxZUZ6ELdRePhUiT954RXCCK28zT5imMGZHt+PTc3VT8HLHZqBDFo8PVxYokZMh189xWVp
i6k7RZ6m9yT00PnKAOUYustIU54yll/z8N4b7LijJ3tUkaBzSPy+ylTP4+GvZUnmxKsGqeC2KPvb
UDCjgNO+nX9rdVtiqS7MbNqmMtXzGw5b4zI7cxI4n8XLYF1nXT0aXZhCOE1395aKxeKRqHRLoROV
EvAz0vIsQNwKwkSRF89SxcB9BG/hlLmL2orZzmOJVKzxw0aAD4siEAXOtRNroSU5g1oDNei1NSEt
Zg4yafP2XJW8z1GpiQ86847ValnON9Z3tqczkSSAQddDAzWo5XVhyHu5mwa7jQtIk61C6hKoptbc
ETIm7IGbYx227UvUz943/qZipIx0MzllzIJP7CRyk8r0CLh96iFXetJAl6O5jg9RBGk29byY9Nt/
7ZyZWXcuILDsVpSlYK9RpyipRL3gzSb+AkZpF5XG7eSkqu0743/XBZ09rbYTIE7O0HQNXZxlmLSC
ErmRjGBmtuKUSpDKRT36OEkYB9uyeB9vrfmeIxrdEuCCOMvbgXS6GwEMLjGLEb5dtrFK/bwXkVyz
yAJ0EFqlf16Lh8S0C07CovIEQNjYWT8fLpvZT9ULpDeDXsS9qrv5U33M8RvuJSBy0RCVpqACMucX
iLg50rnV4ofSLJWQ4Ly0Ec0PxfESQvAV7Aghfsd3DmEqloH16geIfAXngsaX/JZr3WXfy7LtfKyF
iFWUcPWYh/YWDKA8TmhIFkvXvSAcW91bYzFwcWBY0ZomURetdbbDX+uy1kZPfSbpedtb50ZXi1xL
//Jm+czKSC1etZ+3zSMndIw9Fa2j/kFo4bEOqhTFY5ZliFBUQTKm9RbqNRArh2CapIpumzgfKuBn
w1EMD/qPJHL2FRP/MccaK5Icq8rZeoC3n4X4Uvf/8FyrUuK61hT9QGio/tYJT7HRtfJAk0Z34tng
xrsF1HF3zABLFWC6NM8Vc90m+/Gre5oZglqXFlVW3dsotuFPq8EKRPOrWTM/qSJcB+ksptP3WmS8
R6BCCsJ4xIWHBvOMIIySOYE0hLsc3Qbj9uwmvEAwdXXxLiYm6VRlDQJqbyAjYtKdyBvzoKYb5587
S5Mrf3bAxJF5HbZAQKdnJjWlDiYveqXJCWuHJ+h3V8sw687lvLossRliSuVjPHQk8r6hVF6XYJBP
kHuHm6EwkK9i+yuSLi/dwR8DCu+BEOX2hB9Y/A8G97CgGjPGEXE1lIwOIIQuKx/CU5aLdsEO6V3b
gI3xTacPzF5/F5Se8CEsntxjafyLeZqa76yh7EgGz5Exe3A895PZzPx5iiuI2ESmhIFqk0yJ7HkB
pfYfTpI9m+uGV4teGL+qpLuwmBvKm6WH+tZojOqjNSm366hj9c1/C2EOFJRkMmIyOLp8OaG7gQmp
THC5QODQu3hSnEOxcrMB9FnUdxyWW9QW8PyMMFYdazBRB3Pl3dK/aqLLOW791iS00M4r2rgZwn8J
zgmhPm7ikWsdElfqKSM3yYL0jCJVzpt5Rqt6cJ/uU0VyVIl16vQq04Ccy5a54V6zo3p+xnOWEHOk
zXxBo5jEPQSwC8MBtxa7wnVVcIdrLIrLS0tPg7Lv7lWfmXe3xzlFeJAQokH2LR3LqVhJGKWaNqpR
ROAWA/BCWmGjus1luSTK4f8AjX8APYiCe3bC7pHXwRuaTxzMrrgt8q6NPoyehKTD/vOOqgaRLw+5
1VHyhx+UDv2ImqejjCP5YBiHk8AHSB+tCD81upcTavY3ydQtVkfD8esG0pWClUOmrzWtIxzCpZJP
7Rbr7nt3DSk7NV2Iwt7pEEKQbzesraG400oDdFgTa05avR/9jsOxEXlgudSkc5lb2jqY7Mv/jmls
KHLA2GnUhxeV3505Hq22a8Aa5LjLqaJ3U2Ygdkz1231LYHvrTsrjIEuWdtJtx2RGyvjCtlDXuNYV
yA8xD0W47AxaIheuwzVFY1CJ7ARM0YQJnxX97Ax4EmDPZhyhoemen/X7qKyToLc2VtP/DK63voLt
8J6+p22amQTy5uIVeAju2DKqQ1nF9h4MNjWpaWlV6mO+8or149Z4ZVny0w1DlBji2/POPRV66xlF
wC2zew8N4AlvH8vKEozSOFWTasascAKaTvEcEDa5+zhiNQWnZ8WGhkkOQngalKu97ms6GuU08WM9
ROhPfML2CsbSRva2WKkm7xIvonknDkAFUF67bfvcbfwPb4EDor+qsCQup5SveuknQ+YGToQnv0vw
VTf2IStKjTluflchS7182nvLgg4JblIld/jIGCuqRf9ZSsM8m9tCiNZ7kb9gFF5jHBFbOCh0XxWJ
o4XjGMMgRfRkmOWeQ5Pz+O7NhLsX7t8s6NQjJB3UbZ1is4HCv9LmCSLsyHwWksud7xv48TLU0xH2
MUYY1gDqGBRNFJXNMr7C5l8oj3UZ9hvsiop43Ufihpd3ZvYaHtn6w11xVr4ekTms1zMY7DDIIYEo
e1hBnsm8czvmSFxj4x9ZA96WqMI9HR/CpSlpUrfb8lOi4iIJcq0ayO2RM8y333E9WbmShbUFY5z1
8Qph9AcN9ZZ/Ouwyf+JJvXE6xL6CpSGIWfR6N+66SvGz4gmrTG2pe4Sl5gmCp+3sCMl0ic0ltcuZ
xEHBEi/UkPSb19+XABAd5vmSjcNnxNLHTlIO7nMPshRaNOSU/aakl3EeE5vqi0fUkm/GSdNjy2EH
+unW7sLn/NsjJykZlS2JKOsmcqxZJs6K3d6kbls+l30c+4nTzMCB4vXhcvk+o/OiCuYJFyaBUqxL
GX1R3cIzdODqZDLzOvg61umf096zsT1l7B4NNixuD1p+ZG3dWVIpcTBaYOqc+LDk/oNDl1dvE9hI
56hbKbpPzFOAl7cuS8GIJSadS0BrE+41P+xY97tSWjO2k8GXLXwN3gCPQBx7FZgJzF3M7fGwKV25
tJWs56cSYjGzsyUbCxIsZDzaCXLWP11YTZFOHbz4oUTRWbpOrUxLpsvu7QA5mvdnQWSu6savjl6N
cHW1B7r7Rk4vg17fPrswRffJeFsO9mC3jA4ca1hukExsr0F1gFKsWLuxNmeg/z3vYsz4wvUifvlc
2lswGSagahPXuAbrhp9ZCNYKkpf6iHcEVqiCV4rNqBmI0XuEfsSFk5FU5X8CpnGmCXLw8Pj+Wgmv
zZ7At9CfdwXncszTuqDhZJMoxg1FEvkd/4GctLf5R/UUjzgtuIIiWIZzB86+1akajU/KYSXf66Lg
iIrU7FSoaJH8EGG7vNFj0cFBdcT8BwvJwdbU9AEI9nL2aBhWEe7VLjTAfO2vqJvtH4KozyyxkjrH
+UftbuYVOw+QvCOpm/iE8saOaKtGSPfBvA58GGdb6PZc4eK/NvXvFFLl27AAOTNXdH9McpRcO/XS
B9lstb3fud5B2CNVkTBU8g6NGUqluoyFwTf1BDOL3HJ7iHnfb8yJ/j4ylCNPmKtqEZNugMlYjsQE
TPXg/S+Ii/6jLSrZfkHS4HKO/Sd+AjoXlzMu/ZS3C2pj7HG3wiXdeQtgBexCyhd0zRKqxONO3528
wbwPHUK4uekgN5Rs18Y+bZC2ZGbJ9+m40jxIy9uhllDvylws8fIhDtNhefoqBI4E8ockKlro5euz
T0gA/rw2ekYN4cJ4PlvBGKS2ue2/V827UBXWR96fHdVbBZUDEmHybSkElKzSqTBOYnieWM5OSfXO
7ZpKrK69aXWMCWhjh6G+YFsmepyarApSwCYXL81I78QF6P/GUTMEXWC8TFOIfi6vO6tcaaf6xOFc
ar4i7LReLmFngyGLjuni56UiqkdS4K5FSgyGmPXjlKUw8w+zxu5vdTBl6vjVo4TzUmOuyTHsEztA
/zDWzDginuvV6BxOHjFyDfs0LavkLStL4OIUBCjGd8UvLIWVapKvpnSLseGZFroVgpkzb+gsw7md
LaxYsnXiFOgD8YeYExQD4r7p24+ThfPcHXBsdfAelPn0w9oK4pQTykdofA46aJM0EnuJr0sSDxFg
t894bVRq2Z1aF45soWFaelcyn3Hrg0s0+/c936X/DUe8U2qXiQdbkIY720sho3jmU+mge0cnv8Aq
U7ESwXRQiMlw1TXcNzb4MIPFvyIREu08g/g8OFdLIl1j4D6OjWjuz6bnbiPwzrExqkRANNcl6i+F
A2gJKNKkCtebP3E093UpiKLl8ibAkGzBYPCATIVk4ZvWKk7VUBF4WQO1wPRfPtatK95o/Ccu+O+K
IScU3E+v8x9tVbnztAkCztNQHkGC0HiWfI7Ak0Sno476DaneIR3+knMqTkjxGOznaIzDKayZ9lbN
RdhtdB4dYAFggO8VevhNrdOBflWhZzStieIH+TUdtRGIglWoFxg/nLFB7TYASeMouR2Drhsa6Phu
xb0aIEohrQQM7oyefNZry/3S8PNvJ3qiwSbjXECH/PfLtzfHAuZWu2iQMN4kGlYRXfY/trJ8/2Xb
d2vfu+IBqEbLJlVV0q6x1aXnBsVDzICTEMRFySEX3uTS7W396ALOJdzg7yRJJ3/+1uwziGx1wBhY
33u4DtGy5YLhDC7wDW8KiL+W5d5rn7OMOXXrXY1YvPGNQuOXe7eXE6RSfpmdIk4aNkoYSCAtNQpm
ONb6G0dlbN9OBNBGdLT32N3kaGN4yiLKc4dIvF8XTUt5Wxd20vlFBiFJ6s2UlrYd852AGxJ80Ytw
JreKnSYXb+LOzY0pme5C/igdcuvAKxgL1AyN6ud77BxnmSbiu3B8J1aJnQ9xBO2l7kg17/eWzRRu
UCZbGIazh6KQEA296Vx6afCLwpjj8hZKeB4RnBFae93lFTZBL45uAp09bGO7qCIj55zIOx9iNFa1
uSvZa9k2pIL7/3jH8HWj6kGz0O3orT2Y77+F+zzO18TUXPBves4Zkk5kKCp5Kn2vh9av1ZH6TxeO
f9xRP7wpDNOrFsKKKEzqUkqtL5Z78zdlkcD9gUMvIVa9MkHYu7uqzOdLqlOFiJq+BNBe+ImO8mwC
m0MAKlR4FwFE+WYA6WxsWgMkMciR768ywGrCfHzIFW7N/EZW5kOz2JRlWl5A27o4xfSleLz4Zmn0
M/gSOAVGBm4ER/huy0fr6wjKLwI9humDJ9mZR2s6k/GxuIXexSNNe/Nkp2D/qt4CCzYz91HRYvsB
v+B25CsfddaeLytWVEl7b2fAqo9IRQj161F7v5Jpds4axT63R/sq4TTkXFZIlrOiDNQl1XwM4lz8
FQzIqrzm/TaCoMmQ4yLqj7r1zpVtCDGJ9p+HgvF4urPXORLkE2m7P/0sQbe7cmY32bdBFbROrdBD
0kkyUbNdoXPc9eG4LEzJ0REc+U/YAh9yJ5YywRb/GOtBiBPBhl/Ws0q/u53+jBNKWlC6PUR3kTUH
ilSc5zlx3GGRvjvMSv88HhOih8CK+DH9vqBTWXm+XlxJIZwAosBcz8H2hH1MsBJGmJHrUL2iZpR+
WZ4TcmINm6ZVfFjDBSdMJgTRTPBSy+My5M2f7i1CbyJO/5jWurAUvVhkxT2eq7OpUc9cU/Y2E/x7
F9rF16ECOXj7IiyIM9GXULJvVt0GaK5fsIq5x3d4tRNenEba2/hTxvxi2ocozQczg2kgNURooi+K
mPdZz8PtL+qqzrN+S43pOJjb6fAZEflFEEK/M8JYgPm0sSEESnx/9+U0K6+NSWAYzYa3QNCGii8B
EuKUuTnmNDzZauSkZaRN22c72UM8Gz/b+CmGtbdwyxuKZhe9oavLbtQxvQ1tdKxRpUWtMr329UGL
Bfi9auKBDHZB9SbQxJh056k+rmonrUqslbr8qCCeBa0loN1VVBnmNgVC+jAL1xX32o5q3hcimuUo
r9Mxd+4DSqzT+byHE5fphPFLcPzQTk5EaeRnBbeFYzHrYr/WmafVTlTDVWgghkYKTkW2SC5lWrh9
pgYEQBPB+rC2gGby0W7bb/l2j4eZaJS86hioCxGMPF3pm61mdmPOUYnmJcY1GKiRuzcvuRj4mRJa
bH5kqnbBDOUsFDYC1rPMP+4rnEI7MwQxh6ZHups9ZEAWmrLmojyBTAuNsQSaW5M/0pirx9/NFkxm
i9uWv8+Tje3gGl6PkUb8EcVDmICNI8IoshzdlXiEukgqJSyA2ty3ycVogHDOJG2e0l2MbTzN9jvd
72zq8MUL2oLXHtfr4B8nyG88rxDZXOzsMqFe0t6seWeoPdyU4tPndevArYLREOLllg2f0mq35gmQ
syJ1Z3v1+JaeeEA29eXF5FKM1llO/N3w6X2BCcy4FAuceC/d/yQfGDI+KBZF+/apssVJy6b5VS86
1FQb8o2fkg2qcbLm42GVT227GlsIAEjLKwfO9cm9uB05HOcz6+3tuZONvImbZBx2+iHBwSP0MSCL
6APJVNG3FkxgaIe/hRX7xCjyiS9ILNCBz/NqBzFiexCiKpJdlCmPRSpz/i1LrLtNw8+Qw69CNeKw
ctsa32XG1NZB/8zXG7YO0XvmEKvaecJgCx5TCQlDKNvHKsPlV0HUYN8HuCHlp0Yjn7ixRLyjqIwc
9qJhHI+5rYBLeo8iu7u9n+n/AYEG8QgQ0ZsiwDa2fipDReUDVfDuXARz6ECZ6BQv6dvqRfQASCJO
QabLng2yHsN+xOiH8C0PrqLmD/N7N8CYY3Zd9vQqPNJAQM3Ptcvo5fAyr+Dp33WTPmmiXcXMb6i/
SELyHN6SzxBQOvmMmhba/j5kD0nLhWRUI3PWCpVOro0j+DV7RHR5xvsIRHivAbY2FrnSdBa389AQ
GI/2O1c9yvwkIwlx6duI8e4unDZKzFupnKGSOUZB10MSI6TkasG8RiAfQ4nCiguZH47KG2H5FrOQ
tkKGqmFlMK9wZBkh5EYBaJfdrcZPuKz+l/yhU3RsJzalzUGrlkyE714/onr4E7DKIr2S+pQQXfqK
718MbZfExEUqEPJJIDoi3sINUxlnYE5hw3rh3x5dgHrYI4qA2ci9xl4+YsulpS6l/cHYDvK6rk7I
ZSHkLexXPSnhtlRGwR7FEXZMSxaFFfSr5rnmanaRQsCKgb1McbFH5dfJhtKJDr/T2vt32dfh6N+w
8XXEC0HCtJfJEDzVKPFppGk4PhyDQZCXDeiO/pxQTby+cwzFJE5qokdsyaTidYGwFTFbqxI2npbc
fOoiJvV7jSIjri4Dql8RJ5TRHzpzIMIi8uiX+Xi+5TFE7hm5XvNlFSbPhlnzESbTUAYLMjq+zonX
+r+kjk5roaj+5GQSZOkmIuw+D5DI7Kd2wcYnNrXt+lnINNc3GxRgC49+YdfEtAc3PG1dOtKQyHkN
OzTnX99BN/ZeFr0FIyUXnFjKAk8QtIZ1OkERKpuHMyntcBCCqTa2q8h7FTHtuImRShUhRAGs2y2v
Q+5RpCUb5qDLF9kMlpoXiCoc8JbpWl43iRPwEQJ/z0ziiuEcQrCrukl2FBJ2k3UMRnfVi/3l6J0e
J7/UX5/eeeTUwOT3ynsnGyhV3ltGWaDYAwfTk1zNSCoH5MZNdl2+CQJ9S87IPKUY+16szLNOtrA3
n0UQgiinaCCuXt5PIONR6qI9zAKVIMb4yY7Xu4idV4E9yU63DXeMdbPXNtxX+3UlxwFdbm3NDul6
9NZqbxpywAfaeFPo6NL8EKfeIf5a6ZTRNGsEcNsLtBDf14Hy0TkdKcz4eJOEKWPDGYamQIJmVHFd
Zl86L8vMfJ7Ik4Bd4dB86gdIj4ifo4gk6wX7pmjHF17f20Lg4MmBwDdSUAhAA9ZZz3GxOiUHJyHs
o3b83EYLM3/4nWcKaUb4jeMgeAj53YRqL4fqoPztk66xbhKYzV9Q6FgE2jfDLzMjCiW9DCBL9Gqy
nnNh+6BoDSGYwiqqcU7LOF5xKTCBl+j9IB13pjCbKi6xAP8nqcy3z+s0r8QNsqyx3QmUYQMqYxYA
VQtzOC4jaiX5vF2usrjR2xcMLH7dwdxKH5yV2Fr3+EIw7ik+j81sWL+4yQJpyTxgse7x8iMS+q3t
eZZeMVOz32Ml+Ix1xZjKbMXH3LBy5HUe8c8YgpD5YFl04WcFUE4uXCBlc/hvkaWZZPrRM9L9XP+n
dLaz7Dwh+h5FeltXWzpOU9TfjRhbjuz6uBj0iPaivPle2rLuVwsqwh4jHFJNs8Q6VsJGQwuB14Tw
U5odIUwpmTRUiXfazpjhZcHM/NtJX/uqTiLiWmP4pF7QJs2SD9jSnMEHei3zbsfXISJ9vHTIzpW+
zqZ709MDiDVspL0efBbdVeWQ2Yv9DNtFCEUbWn08Le5fvZl3MZrqYWvmcq2KBvMROdBWZ61x/a1i
Fsjt5LyhfYYPfYqJ2OnHw9QKMtj9FIAeK3vMkVsaKYSlchlXPiXaVIrUeUObwCCmm/hbNQZr80tk
dOg5KJbxtlRwamLZJagyVp6eQuF2CaIaPZVdMmghf1ii3V39OsOxfhH4Q6xhaz/PELJZtf6kSTyh
JkkLb0Z75nbphvcw4Wh+kvvHefv7DAYJgqxfmz/qsoBTtZqsZauUHtvi6YgDXmWYza3eMoHU+u1w
lJW1O/rUF+T+Guo10h38CZotg5BlMgfPd2bJW5H9qcVM6ZWjA+UqIZigNGnbTtFzoBek9se0ikSB
XKJWDPc+hjAa4CRSLGHe6ZVxO5oo4IZDuPrcA/zwwSm7MCRwuPZkraeDSIsPdAqMvEhIAdShokRI
NPP8q49XZDctYunvavfSEoDEOjxGeYnGk9ZN+N5el7qbil3eyrUGHDJrxdhpbfWuGs5vrwhqT4uz
SgwqMXVi/CWKbeVH3PfGFt5CzqQXEJ06PJfBjaUTg5OET6fEXKQePvbNA/0tNbdiun2Ua+6Jchrj
ZUHFfrl5QI5jKih6wFfsjG/s5UJiOBDHs143qwIQc76QzAyd91QKRn+Vx9ebV1LfwNEwvlT/7QHU
6KM2RARtuSueEr+7Y8zPyvtqLaq8VMljL/oOYXydN5a3HjaYkPKs3FS4jgSs6sxYk/slkkikhicb
9vSbNN0bZ78NsVrNJ02o33zOvukI1be+YLLZgwCv0PllfuEEObO7vYS7xKeQb+aIEk3JOuIUn8Ta
G8tKg0+rOAe51aM85r7XS+QBGQkzPzumxGCsTvsBkMXW5XF5Ir/87MhpKo+OxboYUcs9uYrRPWX5
ER0R7mWCLYTqeM4J4yAXruoW6HLq3TxCT4/hCSDWcmRYLDbb+6+arQTeSunNVnFKMzFxyxzZuoQP
g7nuL8kMaxh3mUpc12+NPQYcFLOBgup+5JdJBomF3Sa/eXC1zBA6RY4ZpxrKDs/qVLWCJRloAdkd
wNS/gskb/EXs388LspcHNhwlHdoLr5HVQS+nlR9KViM999W8ymLDDikK88YOFrk5K+X3k4tf8+KO
blipL9UM6Ad8bA/9fe43Hyo4Zn4V0+MEPMsehiyS0TvGmHSXzu3esP387dXRz2A5E6rsY+j63anu
HcN1u2abz3acVeEAL7klAEIpufMX83MT8i2/WHmR7FkbjH4XDs88bA27IjTj4cFsIhRd9n327Gw0
V38+1n8RmePvbbZId5tomcW8NjCAY0VX7uE1Bvm1NPF0tUNx65zRSymmG4ZWasHPgQzpnvLho64l
QRDHs84vulIaoYqVm4oSeY/ad4BwzZZqZV/ov5j+fMJ8OQX4sIA6FH2cPF6eAScFMnsspOJFmIWL
/Qy0Mb4QHndpgwpQR8d/Ep+Db22KN4I0cTdow1GkIJsX/oI8uXT0jeIsGKz6H4wjLWKeGuW4LMvd
X6IctSIFhWKo6PuWka3Epv0Ta+k07Y10+f+6G3ZnfLbLxI+S/kR0n3rXYcwEp7k9tUFAuZb0BUJv
0girmp0SlnsFjn0q/UiijaBoZUXVIHAD+PjM/UZQ/5VX+NA11ZjY6ATidZXA3nNs2dcK/IsPhwWa
xybfx8HQxhgFVsOlQSmgeFP7U0KcAnvaJqH4R/B5dnB1qxXqATR26gA9L7wzQGFEfXihfrXyWw1d
CxlUU4Q0pJTlO1ezB/0FF/vBJpQv4K/KYLWMIGuzNPqVFs8QnqLY/WB1qigWSmt9v7yWfdP9xNPl
YUdhQMC4kuIcNGNUFnZycUQxYIMkbUL4ImOaGR0oD112w0lQ48FlmfO/92TjE7tKtxOgl53FkzOi
VlsXfEU1irDrf7t13SX8D3b8lG8H2IHenjqf+iCxx6EVCW6JrX0YCCLOgB3J5X2hH8ELOVZz1mGS
SK62LMvg+xkQjO5GZvH7UTgrfNrdkhgOsaXv8UHZ8F7AcoAYb2mczWUc5rDj/tKDG//B6V+xaNqP
IGr6WE9HZ9ndfH0d4iLUa1Y02+6MvcVZkMBD3tqFw6O9ehMJq7sZl11rV0H4ADxtC3ladk6T5pGx
6rfTCvaCYXqtHBL00jgyQhReDhM/JI2R71cruM7q0n0ZeE6EuiSLpDKh6fGGxXOahnS3/+BE4rO7
EWcpyZwQa9DDEUaEYUsHuswCKwJJsEqpVrVYmA+GzbUMaM+bCKP4MZtJ5INDY/xi1oo4P9CVUnny
73Jcv0Oi3bPhuvsPxC/aQzpOJmoWXe2EiVNAxV/tZKnYK2BneObGtmSehM9QupNWfnf8ycZm3EKr
96KSyjAxqJVHoYghElGoBAkWJn8EISaQpN2uBIv6+m+nNqIKYT6tGYiap+64LFHuKv2WlHWg1k6i
aEat5P9pR8fEGsFs15abIk7ubJtVNZZrLwpmyR/IPMG+c7uyiLBiurY++fyugaAbeTGua6rCS2RT
6VNT/fF0w7sEE79lgrYHwZyYOW3NA+Y8Qzw8KzpCtvUqQTGGpmMT3m/WY86ASjB8x95c8he0uLrH
YjbXS+h9u02x/G3mFR9/O3N3ya9U3uDfpKDm+CexQ+/K/Iz4Zo1G5Y3ToVmaboLDi0OobcLMvYKY
EvJUAlPDj5ku2NevR4MIFjikjComShm0k5/aAPAxY8dt9bF7nt1qxGjYb2J5bIyj8wCsRVgK2LUQ
qt1lGwhx2e/AUlb0924EOJh0syf2l64bZdu0ksQKFjPZyQ+mlwYHYvjS0IXT1/OqWkMVjn6po8ax
d52BA+QKuwEcItk5uBqCXekfAbK3lOGfdOzYWT74yQ1ZZ2sSaxK4XkOJ9NoGRXTlgeLwu8STu6QQ
RP/xS/10eEzrZfLxRXqUa1j8LiwPnujQqGPqzBS3JvdZGRHa8yFjBrBx7Z/bJNYtaaJhrzP7UJIC
X8UOTsSBdgcB2J8yc3pHbxb6C2gddyMR4MvCQbO4ptZLS3EgFkPmiDVyiinjq7gsuzt4kqWaUnP4
/fjOLF1KjslEYjFAs5nUspWeJ9B3nIWNtDalYiqvZ3i6wHiywGFzMvs73vofKcQQ6VJwz/Su5eh8
6q0y/hBItiech1CQZGoS7l7ZrzfMYNfNIklvpbO3LlneagShZYjCxGZzoW6eakINsg5nwsPiypqt
kn91X04JrQBLErnu8QOKHTFNxoeHeKzi08gQQWZT/KfyzoUoDBf64ZtvMxsKr1vXx0dSMBKgHISW
q/G/M8PV+l4SClj+52uT9LQ6qu7OnFj9csRfgp17iq9s5D8rBVcfYwjyqv3y6p1xUDudypKnOpvF
sldCcLTxQKs4//XmPj10kvRwcouDjprXK494Z8RX2FCgpfxxmX9qO7MZcT+1wmY0ye8dIMvQJqcS
DTyHxohjurJG/hIxrmCGPdz/hE/loKVg+n0qcjkNfHiO6J2V9n5JZBzWswxQsVnZzJ8aG5pPO2JM
Aq8fynrImbJnfAr3yXJHrFfUbDWzligqzmC4Oz4IsoumJ+5XWqaSz1/9p6HP4lY7nE28BQAMGNuN
QMVjG15odAmp6ABWXqsEPdTcUyfx2mHWM+JVCmspDXQFTzjKcQTKuvgdcG9mDwOf64iAca2mtqB9
qF5ScyvgSr4uqJ18V+NJOAwv6NHtGZqTeCr5KBv/F2XXvtffJN/o7rhqQVvIlhk+uhL1LGsK8v2a
zVX5CRh0V+4ky1/X8HPFnxA3tjJHWOIuEm0Sd/pA+WnSftPpKOfNK2wVM8JogFg82VBZKlh7aSQ6
6RwOo6dQfin6awHXQYoJMUc8A3bJwG+N9prPUj6S4obMzDZOnh8J51BC7AwPJAIRyCPA5iwPAZxB
fMaTvo3WvHH+CaA+p7T0SHU8hkhmXn1KJzRFnzA4Z4/Dtk4lYccwGH1D9slRuwYYd2tFCM7t3eXj
FHm4vFmJ7Az6bX1Hy630/Sr3DeHy3bPBmqTphoxyuwayUHk+jPC1Tj+xjiqM+gwLSueixve4A76u
nDq4PCsyimlNEcA3zJ2TgbHtvFVLXkSeKo0CJuwoorwv8Df7PaBx19s6YXpVWa/BMPWnxggDlAyN
9anIZS7hGqAa5+2O3BFF/IKrNMpMZxJ15SaTVUE2hD904P0X6GaLLdYP+q7Rodlc/7OifDClYPwd
5Vl5y++Jb4UVmta2tjJ76b2hWjVdardlR2uwDVBCpi/vR4qkJ8q4qvBkLaZlPFGgppuSjmK93+IE
QFzmRu818Ly2t0c8TjAxcySpYIZQcyVCFN8OinQ60TJp/rIlTvkU7NNxFZEkGsSlKqer+jAd4g2T
dn8HUA2hHDL6cJ1rwI8FY2NW+nJ4YCnSc3Em75agwqYEIocRkN8ZHUWIeAukFs2qTTnaZUka3gug
fSdR3iyVeeUi02TQ3ITtyJ1p6eE612mIxK9yZbj4LmGQfzKzrznDMqxlsAlYVB0CWIk3wkPnUsmf
BcnHhfAEH/+Rjuyskmi6xb6UA56WELTwlMKk35ESu54qVVIdOYiXlqN6CDUrJ7wtzMxYRzuG0iXJ
v+1VyqiIjoS7TylPClWQJgXQ3zbUUy8jjz1cwEaDpMRtgg9Q6ytYHM9AxmgIj6FWLzbV8EDhV2Mu
JMy9FyvdDE5twKmaH8RXkfHq0X3oqLJ53BtQbfnYUIsKaqoNbhlTxHKTkgZvqAnbSMgkA3ufB/Mw
jHk4+9tKmPceZuI8qP4Kbeztg2mpBF44djHysWVGSUPEv6VyDZK4TXKyEr3A83ULIYroJ5hesJyQ
veoJVWsSr7R7Ypu1kLrC6f/TXsLU8EzmZqYlBVg3o1N59pAyJqe3vC6zOLUYWERCAHztpPX1YMKx
x4umULes7me50iTok4bJZgIXiWHAekQSivz/HGWb+RLTZOUfbynUhvgZZQZh/oMyW7OQwb0iBidQ
sHsRkRT+Ylz4b/1viPGQcgTBSe5Db623N1HrgITGpVX1p0Cq9kYWh/1gvWbAFYktKRAD6iRfQLeg
FVG3IIdC2hJhxkhoCPI2w87XZr0QxtOtRBtYLGSAtKaLVS4u5ZZyl+IXjlSBqOURyF93tGYz8+mb
D3YyWfUQj3wwMws84xAycPK9M2/6Ys/jQs6LRohw2OSRDZH/AgpER1IUU2LY27ri/D23mu3n0FZR
shQ3TpSMQfssX6VlIQw+cN0yd681Vlr0g5KzicURieD9t91/k79ugaWyyXH3t8oek7QNKie3HdAC
GErX0xOEonaHw5PvHJVGPeZMgkPLhDkERrYQa+mVJISkc4bvJLlXZLzXse+jfRAkVN4rxA7FMjkB
oKsDSXSBS+A4zlwEXMJQt5bRNS9AiN0LJTzj7eKG/unCgy7s8VbHLXIUGXIpEJHmuOdBZNJpvFOK
9mkl//yAl1pZDu2bK34gujuPQcuG8F3oZd0JB2LM0nZGkJhZ/ShU5P6HB0jEAyLUNcVcD8ltsuWp
n7NBOtfmDzFfLHE0nievns172SjfOVlG64Ym3NhkHNX4yQvpvzEqJs4heJkDfx/3/4y+QxZVbbdF
nCzW3L1RyIw0Pzz3dh0nHsY2Z8dzAsTVkRGbAd96iyMabMZcpsbOXe98VASs+93hqsg0c95q/d69
iJLarjYUX55rriYuwliyu9I5P1qxIhAylO9CZd39foqbq309KSpzEjTOkS20mgn7G3USuWW8fOk/
4tlyFqfCYsvGN4adSCUlSqRkkcdBhMArV9/dlksBCf+zVPoFIPyodd8aywF5ZwXGfZbbXJ5SK0oV
kMD+awUHokwlBMHowOw3LAETei56jP0otgkENJriuNZApqjM1TxnfQ3WSXtCdfZH6xvO6n1Eaork
tM/GKgVVq7IUwCJ3C3msWKL1tFpBdM2GOZTDs6ffed2CVK+DTvXWrP0eAs5F9Ao+WvOFvwWq8uVZ
cE2JKJMl843IzUY1460TrvLYCsiXp9omo1bpcB2w/P7+h7JuCJIzd0QMuPylCDkq+CsOvy4tBgEr
y+889Prv/5fV9VxzZ+bKem5CNhhDT3Nj3SyYGSoE62PAgQLTZfH1qx5MixeuLlm3q2bXKXiWW3Cr
ERbrR5MfNL5O9iT53QcAsNfbIQ3B+v0xa+U5t/aBhOr1T5Ioafd21HMvnGE0/vJAQrZc/1teLpF+
P8qYRelxPIkAv0u7HBGx7nkYolGJJY+8SY09JdWx7t8V0172Ozh+vvo9erEOqkzVNRHhK7HldXCr
2r+pNlKJ2/T233Tw+6r2r0KsT/6iup4U5ZisjnMML8KgjTtOozfw9KYMs8HfH6fybzG3oh3B7Fkj
v85MCIRtjWyWxJwdEoHJlc0sxMyIWqPWEm4yyDPMS/CTxhbHDo4F3v+SO6CVY9CE3uAKCkZ5MHAU
wr7QCX/ieWIoArmD/YmT/+EtyUDzEhyCHEOYGCtKXht4jWKCGZL+xPg4fZ8C5bNP+eibbazPyHfW
ipWSWYRWvuXsObaqJIVDeUOB8dwmIh04JYxfseM90FU2EhT00NCHxvystvww7EiyShhuIQHhdQuJ
toSlnfTSXub6GmHc8LtZKUf0MbQhHhLuy7PuhxvF8cc8IESQ587teT48T5LgOZzQyw7WASkXTLUm
M23o8+n+JY836SN098QJ3edSGLYxw5RQ2yiDxnhG8kMopi05x3EzsmOehm2uk1MyUhZ/XfcYPd2n
XQVIyO2muNZZ8P2O60d0oA2Fp5SFDMmhSGYTMPfhiI8L8U7ms7dNAinOKavxZjmZK/6fGgBWhizW
SAhAoTSB8wfxixYe4YUO64za3L5fUmIh2qxEDNOOdMBzSnnNgyA6QpLFCpEbBhv/srEOpWTX2eZF
7A7vwv8VCil3OkRUYlex2WbyejnwxPUKJxysQ9arkJy3uuuT+hjD1dfaKajUcCX9GPZP2H2xqKHa
iX7ucuAE6r3Lj9Zwty8V3jfcgbpDGde7MFmtetEvfgOVjIR6c8/MZU1TucPLdUYTTQA/AdbVkmY0
Uf1NXgySDBakHT2XIvQuzzjvStWBSX/tHg2qFLxPUuZaX+2QFRzCWK1xqi3p/y+bUl7Ppgl1lPQD
d+9JeuYqi/ITLevM6PFDI3L54GDRiJSGyW2vOf3R9xx74chKLIU8oFZpf2caWPkN6GtO60coGCl0
x6CN4KplhkjO0sxhjAIovYWdqWayyGOkIVlDhYTrd2F2jLU7eSBaFxZF9NbRIxMuSwNZX2EqJ1jX
o+mX2WCTAk3dlf4e8DrXqidiUkNGor7Qh6/SGPU9ViwigNWE4msWWnlbFH8HgfHPF3kWsdDoMFOt
/HW4yixP8OoAHMhklGsup3MUvA9snitdFCyXjk+3/cAknKzL7+9nb4Q4XvD3kq5Y0c0HotiUVAtK
q2ophuUxPNUzy7u+cpsWBJ9+s35Yn2ZBHU6LiEVGQWyZcaCLD+m72e6jrxsBCy7aj6symw4iX7ev
qebZQchEheW0JegwVyUnxWw48SgCkAo8BZPZxTUKCbbKHfVTk0reiJNcdPhZCCchUFbS/O2FyDJz
+Se+nZykYT3aWzyCQgDBisFyAcprR6HL0a+SYDO+bBmBh+8HzyLWCXe97dod8YLiKzvwIRl5KwNz
XgXtWSSNU1CHZKJEMHS/G38LuV+2cuG49UhO2TwiQP+k43y5DxWYlp09A2nDmBGfCMG5NkHCPVAs
cRshF8PDYGmGGdw+/DOdzbBBpDaXd/AXuSkFCwXEiik6sUR0ESbz+qEF54sv9MjL5khUXYv0OVgL
b+ScApRa6gPW7iR8Zi+o81V/P8eNlyTRItGpWCyOvUtlrO/jwbUFxj9YlCTC5I9CPEpB1Q68joAA
pFnsncqfpzasUo/7BOC0jMEbG+ydVJqhPnqm3NZMS/x6LausZeLoo7uDQAB1c9NO2nMuOfvLGala
TuX2Y3Jha3clNpTztyEQ9rdDqY7LVVsUNV1wxDO/i6fONklHDYnLEcd54X5UNeIrmSDZ61Wg13d4
pewMGdfITF7OiKCLjMonfIkKKfhsg01qyWzVuRTFTtuY1n/ltxTbEiOLR9n0MIyrPhrlXUmfJvoW
+sCNCXn7CVePYZA928ki07WAsl2+IEsRQ3yYRDc0AlOGDNo4Qu7/QiZtUGk/65owjRQxZd0NRG4X
fdPZv9a9qbDXiaEumHmVE/U+yUlv++ZRNnwjtsQsQP34LmtKZvHe29shuE0QBrp3jcyPEFU9+VnZ
8Uy9LVpdK0lMb8wVCnrraV5OQPDj6z1cLCrleLXCxaizki3mF6xZUxxXMqYSqGnGiAQ84HP/YWKP
DUgI6y8As61XhUJAWX70anBfsqBPGQ0MP6IEa6X7tPFDdzO8rivEeaPTy3InKAn5o/3/eHzsFlpY
orpwW9uDhey6i1ScaOrEYMMDR4MfoDDkARdrTW5O/uOUXPLuVELqWutVWmmvXp96grcGtNQt2rhh
VHKzgUndSWsL3HWRV2AhID1+KntXokIsuObm+9i2Bm9hDFowuZYobBYkXeQpGBmSNDbD23i3qgdS
72mwCP4Krk9NdD8u7c88Da87eMDjGwXSGtMFOxr0JRTuukvZ8yU4e+dBEg3OP9tQDU4m2dLHV6JR
vKHtChHfherUWUF7ci/uevP2Hrb5+HQbUMH+wt2sxELI9dCtgZ4Mqe6RyG3inSA1/W9UFMv4gP6f
bgqZe47hLIhQzcmDxkt43PKO5UpgG9YFBeZFxbqb11ndUuif9/I8B3NHD8Fp0HLG0SG0qAUO9wUY
aybCc76wTEXhU/7wTBLB/e0IHs0aPhC3+fFIgLjg5BP0FFW5Ul72URx8SsjxvOe7Qw1cYJFlUo4L
pfzWn2y4x21QT3Mp0tyxg9lpC8Yi1BZHXMosPfsyqW3CRzA6Kv8enbMydKzzR5YhtMUNKXaSLVlK
dl6LQhf4iW1YugQIgN64Ev/is4aBhWovmXFaMq6MotCXKYE55hxrI7dsckHdkCwEc6v+KoxRHti2
vieihRxur4K0+T0csfYYsXju4+1vknu7dvj1rU8qDesayQRHQJOyMwcbD5lnJlx4RgnysS3X0k1u
mFDsaxc1AJYDQceskmvlNSl0GAyvv0gIc1+DDtBSW09CiNzmfDR/0rp/C5k/Vm3bzt/KNW8tD8l+
bxzWLtheRCxdmDlqLEbCTb1B5JlCF08zMwW2kwc3mB71kjOKsyvWPsDCH3jTfScBqRtj2Kg9vblx
yWinx0j8UmLbxs8C45CT/A51lF89SRrk6UUkCFqPtskwV8YiIzXOqkryqrDj0NpKSSoc9BW3Ye2H
qRYHQQKwTy46bUaOtro8nqCcDLV+QXUyRqcfa/7A7dklXUXVLMvVgr8Rx3wpRe1oI0AqsodPJ2ar
yEmKB62bpEPkLEGBi8VLR/qW+e/RXZH2k5q5+pvdpt7wvVmr+NMBAmDqr6B7oACxiCk+Nw9W6WZj
k30h8GBYiMM+lr14rCb4jMA4pvM+tzH474tssBdtTwkTDVdulMlg6A8WZNMTCneqI0fSo3n4VuSk
PffD+lhdhkLqub8CM5ThEDveajCcTiEO8RX99fTO+AgF0hzX1ZI0U20J0LPHYnt7U2rqasRMilKO
GrZz+eVqKGNhDZL2Vy2cnZLAnWNX632084kH7mQ5K+DkFYRWNVaAzRm6Mg4ppg1NZGifH6fUBQAY
Joi49lJoKb0eU0YkcWHD3W4nYT/J0VoINHQ5EZI1r1uiCGiCS75L/9p0DWCHqrfiXLAIhTozr1uq
MwP2BZavctLl5iopvQNgPwcPNvp6/OWMi8KnLwLAwMehBDiYkPPIbp6kpohOlo2tU1ZImdC7/Y9i
6UdWVElf7J3A3Cp5KY/YfqA54EUSH4MhibIlHQmdfpVbYGw7QuxBKDKSluEAsykZab5T4taHKt5Z
xDC3chGe9eenEryPiZlx4myD5Y8OooHKE1uWwg5hh4cMUerjwdnOjHBVYGaqLfdHBTXNLcR9FpXs
X64aWvQTt0EFY/pj+Ao8Gg4wblXthKe2WX9veR4ckbsGWVNLviuXq4pKTebLr2b1hivW/gDmeDU3
Q1FdiKGtFsaTvY9rVYDJs9ZR7AaJDwvwTzDgyPbk0h0bEkVI3kOGGzl1LWaV/Y12w/rrD9OfEOCb
Tdu2ul4cly308V11PPGa2U25p97fMUwC6t9bG5tU+VdH6VexRTOlD7vEPTQznUDF7gVuj7nnwKiv
X51saS7sr9yFmQjvVslCDt+rKgTZHEhsZjRICEKfifbYj77EN352Sm4mmgzGH6msZLi1cctBDPza
aH4le4Naxk2UUMWTQ8/uAMw5/PEEOLWLnVTPi/HlfxznkaEcFAPyD5UaGM+aTXEqJQ7FYXyAEwq/
9nqbaLEf/cXDodrGsIs6lrI9La1XRA/Zwx+4vSq2Vi6HbGjDBp/8DJqObuby7sgzrI6ynhw9LI6G
IvWNUdIlKZhBm5pBt7AHZgViHsq9Oq5QneDYZzWuQw0Tp77c0uRZEPPZrBWu1Q1Aybo+l/LdmCiX
2h1HXOL0VAnP7io/DaX+adhVJ+mlC4UGGglGTTiqvbjisFrUvHOXfBHyQb0rrTrdZO95pt6FVegY
GDeOUVYuB3sdb/UAVicZNdkX2Ii9p29/dbE1vpT/CI/q6jw+0R9r1AMoaL+8KzBfJLvvhYEkl6RU
/uMe1RPi9utpf8ySaYcxVl9XJ7U6fBtEMFLlwqAEgHsPnmPSU4SowX0m+7Nse5XBuWof/YFN9PVt
SYwFkH152clSo5zjfsbJI+1bHQq9YaHMfCQKBNpT549VikcCExz/p0B2AwT0MdBXP8jqoHAe50U+
yP2CpB0Nc8x6YdJ07Ku+f6sTtuLxP96F/SJ8/qfrK5mMJZm5AKasA3LfIvaOt69D9adHIAZ12Qwi
BIxks/ivWG42kzq88JLI2HArAfMC1DSPL+kCWWGiP2A6Of8o80ijXpGpC+M1XG0ZopujBzWKhmj2
3iUpbvGw7t6DRwwx4QI7rEzQRpm6QDv46EhoP/kHcmqbzKwR4JlzqbwlP0nx6W8mEm7MLdlEAHfV
PbsK2UG7jWOO7ppHU5CCzrVKtK0saRNyjfKHygnr1ONuWmTCtMPvy9JYZY5P3Hg9tIJ18ltUK54s
nx5jqNKhdvnSzgjae6ZbfX7Wpi3Ez1WiHB0QSkI9eH3SglPenczRv4A1R3gF9t6/QtpIoXZboEJA
mIkEuaO7yxpVRCUMIUi7cyPtYDcREEb3QijkGrtXZ9LWmPNs9RfDkmuNlY5kpMfFyDVh5a1pyrrt
FsxWHwvovHIZCUUlrOt6MqWYJJY5oUWKFhgf/egPZQhVnaboZ2lLTjqYDWZjbkdwdmLHfPFSTrYc
5uL6XvMa3WJlbSLzNE8WZqE9VLGu3SInHBNVjc6ej2MFm2yIZsPEaxmOAZyTMpE8b/0BIrLNsFAo
ks9SHASUX2o1c6M7tfFuwArp8/FdlxrxhyBH0Ks9avPgIU66eOpkE0v4uCoDwDrWQW29hOFu9mud
nWftJj9m6/8UdbGfDVpOAgGjPZa1n+HIaYj2QeypTVbKflIEPcs9qMQYjLVtji/FLuJgO6GMGKN9
7192+MzikjJNBm5Or20Wdmt68x0fpItnDj7TNNrz1sTRFkmcaEsqgbES1Oi/ZbNU/WB/J39Mdq0z
U07BttNxtiy53py0JicGn0kreXWy7Rzj1qOu92FaMYOrzQOmndWFFMr/gK57JnYXFeuzOkfV7Uqi
GHPKrfX70BzPpODZMr2p8pJM0uR+PLSPXAnDKF7vqsVKMPrXx38FDyPGr1ei9JOcOr4VIKwv8xDE
LGKhgy9NxAP9urVyLZ2zEQhOHHzYuxio1xslttRO8alfdiAy589l8tor92qejdhrIBv1yqRaTYxh
igicJv7ts2WdF32oUr1vz191adscAryVyvttHES7ZffeLfy4Dwir1+DO6wTcKP6hYhlcwuUrwqn8
CBOuTj4UQbs+4jin6prpc3hPlzktCXsHRInJTdHiQhuRrKO3rfi8/vhenGSzowNOsOI1F8RtDBno
487xxNglBMQtjGaDafDYsAVKNzQpE4O0HZDVQACJ7rsrT76TLtTU8PAoy5Z59cT5EH9Nxi7UXW6w
uwFZXZfF/M2yvbtAhfuMK6MBbmhn8tzMuElWvyirn7A4A8KRZ90F4MuJ2Vez+4v1ozI6sUF+Ylpq
RJMuecQGUVeu95iDCmb2xxtF9kFKFuHpQbomZUDxMFKrxGjD6WUydSjbPRdCihaMXMOch6XmLSBb
61H3d03FUY0q3pVp4n9RhUj4NwfSSkcUsbn5U/nlFDvfK70IDX7RqIOhGuTFxMe2o0xx5gy1pU1x
lhyBzZYsmu/Z2fqDBfMKYNoJPjh8xwSiQcsVGHI7SuD45V7ui6hPIJrP2QjewhDo4zRq7z0GC94+
3MCLolc/aThZn0diS/NQLvDNFFV2GOCP7bQUfJbdWonacYtqtVWVaLWcejB19YQ0rK4utONG+ln0
eAQ860wcxJEplnTt+qhNd/d381VgMpN/6Adgck5qC06B5f78W8SlbyEU2PRs3wJNNicCYYUSE5yy
V6yYhj0DhfRj1oFehqasRPh0+fMwxMyscwjzp0sjc+k/W/U0HRSchqqxWgjkC/NvYL+tUUaZr3BW
4ElBN/+WDbKBBYcuIOuAYf6J6g6jYuKfh8OZaKvV7kVY76ew+yiII0SsOw5FHOg6ogXYBybagRy4
uFYXLyTSkvIBCA0SarpDrHkK3Dz3dRcAUCvz6vM/q2T99WXqt0rAyJi4wo5Lowf1hBoI334tytbO
Ovhhj3M5lVKL9kRF43T+mov0KjikDqkF29NzaMSt4XdMuMR7QFwT8sxtwa7SY287LsNEmCmZGaNu
8msOF0gdMQtA3G+snP96MSUAws4gnt9Xv1oMMRIZ7u5zQwzbTFHlylRWZOqVHb4bKrqzDc0AkHp/
oZ0PqnXIThVcnRugQkLnEgjCaoM4Dwk6cLAszGavCBofzOAPyznPHEHav+DdbVwIlVH0yBNFLPfQ
GH12N4kXekFzPbq0/DvhntgyeqpnGRygTptak+s4qtfpkq2OQnjLL4vnU+sW6+TTnrMP98mqcfsn
w5rNCymr4tZ5PnKbXoe3X6q+1x6787B6b0Bc3FsZwgzsd1zY3JXGJPeS7zbg/FEb7lWMRFiZy8db
TsKfdcsK5sEY+pilC5a5Ms6MC1ZpJCeRU7/wOwPa/9ySheRucL89FkgixoijCfRHVpZW5CABjzWw
+r/lDZZB4eyJ9Y/fD8UdO2XtJcfT/fko6QXgU+T9K8Bc+N0EQZUJ6vmmOj1zGjpEp1W8UvbimRTu
t3QAKIDLRmjGQjx12h9STMQq7PwpLB6U9H2bnC0WzHPiPofgfa+6butsQfs7F7HMqSc6I8+a74P+
TRikiv/iprD1XF88zQmwb90fZ6ewfj6oiM6IAjt/HicE50wtOR5CRpyDZf1ZxDsXziLXpu8qr0Ww
j7HcUN+axEAgs3p8Z32UtabzDnkAkAInCPu6GS3DPIA/YuV1smDaAvN84M7muWSrVD8pKZXW5WVe
NRPmNtO50s3QUwQYrsBqim3a42CaYM/oCTvyX35S0tUbeSGlnhmUgW9KYIG1wGXJEsr++2ufHmt1
6E9VDv/pCbXBOGGS/nNe5TZMMtYvO3zCoSmfEVNckscRGgxYRxFmFftExWGv6C1CdFFxR+zE2Q1t
j1GH/NYiZKcKPPkcT7Bt0licg/MHkrnzt1Fpj/keq1RfkIQN3KsYa8Sq6dMMdNTMmgM6B6WemYXA
mi04HFLTQjOJdeiIx2nxAJuLipi8Sggr4wv5KyKuGb1orx5JMeHE8fEVINpe3KNq7m8WvY+jcfp7
Uul991VqIF6PU31FmVW3oOAiM+pB3zxk3Ut4b7A4EPHJeW6ykExSGoC1DADTfOLo6/mT8PVRxcTL
JM2l7V/UOQPlejNs3J+opA1F6HeZvcbxp1CGn09u9eRl2A3tWfJRijZU7V0GjonIs9RUhOtHZ28U
MG6IoZ9kkogKinUV7mPQiEIE+pggJBF9oEXiRjcjqfDVS+LQtTiwoKPFok6Hf9nkGT9tBnQd4DAB
mv3dM4D3nBoHy1mzrTtRipEbBYpocd3KB8Q=
`pragma protect end_protected

