`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bd0FqTI7c2E3CfpymAa9GMQCAZ3uE3ZypNc6kDliE4knwmFE1bBtuW5m5K1xzhKfnsK0xV84C7kg
8dApxVNEpFDZzInDK/5++FH+3k+QKhSUfWngwBat3p8AyDTMIigB67yTHowVZQhgnXFtwKrH5Ho3
6B+8sqc8RHsCPvn5SCJzbKMO/ofhnkN6MslfM++7oDyV+BTZukILmYN6FAMe3h0DOIibjHvuzgTN
TJeDLcy7zslDrWw5QND14pkFe6zEGbJTuGse1RwDt7ch4bP5PcuQZ79ymlVNOvMVYwbdLrIYABhK
9zAO+JBq9d1wbKZN8dbwm1qlVwUvv1JiyW3sug==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
aEOq+REjbrM6JbyWVXWLCWzNF/5kg/9FCh9Xt575uP4xJANMPGebi59cVejI8oHJYd5CGD5fa0Eb
yN+m7exTlaST5t5L3bAu0Hv4W2/qnQ7ZT+XIIj7XSgmDZO2Sree39jf1ZpDbhVUb7X64Q7DOy28N
bpryF5SJsiJCSr1E3tzlKOeKoXCTfKbt4wMGVhmi5S8zjUnxVn2TdPQpf+Fq91gUatu/4bjo42BU
KHJSd/utVQJx9JWBGyPnL5gAySbiuhUTK34EOfl95PU0kXVFZd9QuAs4YyIZtiWKQ324WmkzrpKz
xfm7H/dmgcMFMJh08Dsjgpn5fnI/G5pauqS0RwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FQ4yWqC6txxIXn6ZHntDzV1u2zLPnlAsS2FJQ7jDOc4Y26mPvymPYNF2awArLPTK+ikIisU2Z7gG
va1uz0VZvg==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
JH3DYi1Y1o+Z48G08Odzz+AUXAMYj0MVbw8dTn7C1EAsXSsoQ6APdZjCch/55LzyxOJnyMEcX3q9
CkOleCK6DqhAqYfoyajKOxrkCo55AFPvHkW/08IFmEWZSO7pt87XHe/Pr1viS3WD7JMptgnovz8k
aKdfaVSzfEBF1Si3944sFcKzTtQZzFHSPuhaK2Mk3Pjywd9uqMVmXrXr7Ponc5rh/Hkals0qVnmQ
4vA3rhForQz9GAgRYH75pkMRh27JcwT+Y5Cx3S+nZfJXgjcPLx4Yhw8Wwc5xxzi/J69Ie+H6hB0R
9qTdYYLE8jmTPYlOL4k0O6Km/XDyG/QMkTmSJA==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
j5pCgBZT3JqKncqbIIHsQx58tHzAQ0EUBB/965i5TVtyaZoU5/Lw5nMBlpNoVE1AeT0wRSbaBunq
YPaMBfigJlCdO4TB7f7q0X4tH7Us80UtQlyABlfnB1EAhZO4fG/urM52tqw5JJHkRewNA6StAtLc
d0DUa7TeSxrPh/CvfPsl+NHnhiVPM2TTnFiUyO2PHLqJKzBz2kZsL0tGAHQCBbi+xYGcZRk0k7wU
XNoF9+KWqg41MPkGr6V9rCXvWALnbO/3IqIKGFoVTepsq3q8lWEX3wIUEuvhIZ/crzMIWGos0CPw
KVvIXhd25WTg0KZw7fC8eXFiVanX+Xn11t+amg==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Bz87fD0+T5j7GN0IlJxgIC0yVYhiLCb3T5J17Sg5336ETOD2OlJU5kwAtnLmrDuTzQ76pJLZe3WA
bAZ9icjTO5U/0/orU8PGzhokY1d80QZG+0iD5bp9xZcqwwKLBDVpgVnSa9G5Dz13sRGxNrn+htw+
wyAAQVXS4iKbWDIocpM=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ef3GFNEr0AIIdyWT9nbMtSA1oYb6sNF8fLXcjl1IaBtasntSLfUdEQtYlTUhVmhJPOQia+wCW0M2
tmkE+BRScrDsvvPQ1biPyilzfwBbSx/ep67FeciphJH8gmksaKeWmjDq+3tePsHA23rp2k3tnQ8s
bnn1ahRiT7YIdSDUL9feHZQu28pr607JBaPY2H22pi2bVRCuhK16KJY8+KnZQsRIV3BenC/R3eXK
JR+KBTiNFyiJ8/2ihkYaE5ibCoWgksFmPk7zhw/Nb0IWunI7Zwkd7IsJ7j4mxqUzxBYMDkBoVA5a
/M5ZN0C7J9+ugzMgsuk97QpUztRDu4x5ZPE5tw==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Bh69UHmwfAHdWp0ZTfj2WpG6ao2cIO+nran8sFOvD3W3Vu88lEpPHJJGfmtJLUkk8DHscbV82wCM
0rK2kTWHWMziuSda78bq9o0I2piXldMCR6tsa+GYVjWnkG9LX5cvNRGLJ4d6XiJFfQUiCGQJu7kS
ueUMjiXDkYTFYNtWo2BvStIg+WGUV8+b4NUIpH1wDsU1coYHUwMRebGn8xuyjxdba9IUj5tOYHe/
xcDpYB7GHkxldxUndubcyXAj1rzCaUFnxPv+Of+B0nVrIQ+vf1zY2S0UfDyXDTHkoQv1VtJOH2o4
M5rtQYBwgVuGLi4SYcUW4/f0gdyAeYIy65IN/A==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
JuxcxeTPJpu6MhSHPn58M50yK+ApufgxPY3QzQ3dJi6sWwesoSpJ6HhANyB5/ZA7o6lndY6EeoGp
qTApvcX5cMz/1qlFTES2tCarISVs+Z1m/0uvn0MpivFKdSGC6NB2fUeYQ06eJlJSyP88jvXw//5F
ZZ9xRTx8JDLPM3bYWAg=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
GbLh+9rhaMbp/FWiYrWxv7J+75aaJLRPTfkykskOccDDkNSO0PSKWBh3CmVQ8j/OYHHDYVARWFq6
BBeVyEZqBLsonameDtpva3RVWLfu8cDDJT/BBKWLy3Pv7UlpJfbhb3c77lcmukdaq+pLmsEASAMl
1XaWO0yJDk10qn8Xx5T7L3GdL7FnKbD1wDjXqZwYGQXsNpdAcbPyZeUY6GNZn3LeE6LqXTKl54Ed
xDUydkpgg0sBnU6vZ3qkNjHQktpQD0k4Igylj1nTSY2RiBz1UeUg0VcQwA0yB88cF9BGw6MO5PfX
VQaaJ8BeW9h+P+FFkkmKYSwvJQw1SGVaRr98xw==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10384)
`pragma protect data_block
4TpDwhbp8vrcxgHFn5qXXuRXxm0E+hfTA2mIqdeNj6fBSppEV9520u8fwBjwEpQvLw8nJUBl1p7a
h4GQcPDB1GbcJgqNyukp6h03Gt1IM5hxpnu4UxDkXGW6CViPCWdJw6TGoFVZ4DQachG71WauJQ8o
lhsc//7ssbwvtpIDK1fGUwL3lrd4yhNS5G1rZFpLYkW/LHtI1i5ZWHBJVU9ZUJZRMTcGrxGSzcjQ
ddMfuptr4ZZwUBs39jUbtUtyDd5RBqvcuRf1/IgCQyLR6J99pUew5J/xLD68z0lbaRTK3/AcLH4K
5KkRiy/24+sJlOCtmj691UK12RChpR+lTFmhtJBDuzoanx2vcJUiteoQM5IMerXVF2R91+XE0JAC
NS5MmzdIcVfhZUZec2mi700SBl86haUUwYdIO2VQnrpPzGCXnsKdCAFeAM2A+q+5aVjyDQFeFyYE
wHvWAx6+XDDgziafMAYWq7txLajQ6Q6H8yVwP1+H0aYtcX/Qv+7qlTlQJVzWZw536fnxRQmy0cfY
evNqJX4w1+zWj0n5rgawPoEZwRGE5JouPzTAD7SMKNLI+w22uU1FeYb3uDtePSIHJwQdy3m6D28/
bv0m/ZFnJQ8wvacZspr3NvdSr/agd3tfDfQzmRQkuMWfhtGlfIar5tZMo2vPeeBLoF+mmjPX4oN2
jGszB8iA+dMbD+HiGKH6/5EwC1GlN7TYI84S89sXfzykI9g3dNoLwMHaJuQa5wrrnuS/A24ibvAO
918yBPajBYOAjDt0yYrSw4GF6dPWyredKhjgK/s77F2NBC/zmj67T1d69VP9d0C3zB6U6X0RUBSq
Rc45ID3K14zd+bIn6Zfih1GiIAuWciCWlu4lt1qO3IUl2H2Re+jW68jtcqYZwQK9mk4Aa1/8Msca
C1KuXgzelZ4bGoPSQrapkKpMEuCEjU8ZylFUwECSQt/4R9TTpMIa19+5uRF5lzutId/tZ0SLCV0b
bxAgSPQ30hPHYN6RJcaEPZy7BnqVOix9Ft62cysQhg4WROpVFpCpbDNxapGxesdYQgyX/lAcu8jX
9OTR5FjRWsSPPO+/XsjEjxc6uVdGEg/56JdxOzoG/ElT/TtGJaQFHwfdl6NnWMnjr7gCgitss1Ns
1p9ggDZsaNi5Xf/SIwC962tIsmyLmC/QCUL2F5BSRbXc2cAfN+wiRqAhYdl2JTAF8M4pAfaidXK6
F0XqcWYUud6voJlUgZ7pgbyK7o4mkGGUoQTvVLK7Ya99AKv3fIrePP6vzMynshg49jPCi5KCoDCR
eSRhwONcpicOoZk4Q+Y11UPsQXbHltKmBpghqO6C0RkxW/Ukoh4GJ+ItQx15QHzkldwSATvIp3C8
2ENnvaE5iv38sFNSQXfkZwzPsRZ8FaL0+mdtNuyORuH7Zl3NqnXFQ8xAamWdgmYhDi7k3hgQOVdn
qNQcwAIxmRCj2fVWiL6YwYaLZbZdb1baB/d5fCiYyZ2DfaWY6JIguJkjt7EoNK9JO8yIfZ9EmGuA
v3SEAhPF4BWeaVd4YB19QjIJSMO/zydPcz5abMSiLZg+FGAHkDYObtWhmEfTSDLJwrtC71I+Wcnc
/pS5/44HQJAuVhD1l2RPJDyRF6rBDT2Q722cIB4P80E4Q+gc7W6cM9V0oCtclRYlRMM7V9kALfQA
x/YdyBojvY9HF6sSTNXYPJdekBA0A/OL1nekhUfq1YlrkyRlkTvrXX5VZC9xzXiC6aeGUpCkrN7g
XkY8i2HklEeyTS8yMO2Dsu4N8OwwIoEcn//2CevmyYtmaknWq4NJfauvWCXQhXMuahH/9cZO4v4p
lZw/E75H06LdYnY6lF+/ok/+4fFAR77j76AkRygX7uaAjWiTplNPKg/CQYEBLJdcrV5/EX3H7r5B
JcpVdCn1ekbXZe+dUSKfill2vPWENY/eqztUjwPYoZ7O1+Hgw0uq+YzOfERBfqv0Y6dair3qiMGD
Z0qXowxeXdYNzszkg+Nzs8/ELmS+PAAcD3J/QPMm7Vu39p7A+7PRkTXbdjOy+zXpxEtg6hnx8b6B
7AY6NPlAiRiRNuDbPNvzde4EdE7qzyUSYrBzucFUoqJTVb7SsweXBWt78jVDpLgfWNqG1tvLElEB
e/JwvwK6gjODk2JcshkDDSozPxJl2ZP7SVvQSA1c2JKXsV4Qxvo9EPZNKFOcBCRex8EMNKKdqPPa
9zRyNMWshxQ4kAT7IxWQBsjOsPomieu3bMEW3v6Q3kRDnwhcwDowuwwqsVEMLiCGILVO5MOxhzKu
Ww7zOhnTUdMdFKZxGZ0vZuk74nlSOxQxn4CK+fL+kGt9SzCbKx5T5aAIw4T/Bee6+zHd+lALqqVf
vJGeXy4U0FEHIDVBT5YVfIFPEV6qxhom2ivs8iE05Mc/oh5SSVTAGVB1rhMT2wJnl29BL35a7336
q4w1YtUXFgouL21csarKA+4YZCyMnZe2Xjg3QtM9blP5l2BsLIfyjTgC50ACv6e1LrG+pWo7LSLF
fqGOeJPvMDMQsGrKPBG9o6MsmsnUnAQXLofr3QN+0t0PP5BwRnNtGY5L7q+EgzXwm3gcr7Oow7tN
ZdJin7fUjXvBqxo0lh1TLGeWZCdoePBrgWFSgNziqoNW5iBmGq2E3bEaKHg1jB7IY9wTkN5p7ANu
QdNg95l5qAyrWYXjWWduklXsbkIjXFFOqSjRjrfFDVp6IyCXhhB7DLYfO5SWJ6ThgchQU6BP/jCS
HrMkAbXRbSyuICp1+M0qiG5VED3hsrJ5J/2oLGPaZgH7TTdXIJkzlU4lzI/F2dvKbfZ5N7SeugO6
AJOXP6sLduPLMXgU9ACl7QwCxYf1sFX86nK8NQXJmYwFsecvscsBaDBjmeBeNzX4XvDvohPg2q1S
ceqi3ED6wgY7KJl18HgUlBgadAvMlzQ3CmrM5s84C2Dl0ajArWiPihwskga2OdFnBMf8lbBE8/1U
z+nHb6qgT4+i5KHEZkvbopfCngYhqEO2XcuxaB9XG8NXD1v1RY01pRJoyDy59ryR1M3jUvmuvKlM
361rzEwVeZpI0eVusYHDHWmlqCYxwoSDmcO4Q7meAeivm78JWRunBPoT7i92fQXEPClOQm/xDrgq
fY9WR+4DFYI4w4fCrvRnpinohE0k37gqO4TTwG5Op5vnatlmviACufS6EQuJE5h+OnrabOBifkf8
MK8oSGuaYZsg3e1OknheyIvO4eLZ6OjOxyXflI2XdKHm279c8ifPzZAp/RmgjAjU843GnmbnDkI4
WbpZmvdbNa16F9Um45maC7FF3R1f7cXXZNDg3NMSZ4C44E9OHHlzmp0TUzDTXD5cWYOyb9KvWSq6
G2wP0+90IjqSNRSQVaVqEUJ6VkIjhidPcvxj2XMbSONupaji9/CYro7RJ9BwyLDULEdFmd+/MDdh
fuzkONDyMysbpPNFgbm3ICUNWslHrAIfcdDJ7wnewtci2OXz08WMqp98/GNaWq5sayDrJHKOmeCy
QHJWeM0QIEMl1kbeeSqk+iUMLEF13dUicyXaAZWgTKNx7KSQGuWB5kZeBcplo5Rnua5mBI2Zxik6
b1xUdpwDiAs1luQBZt6LwG020Az/EitHpzij77kMwc6wTzrYamo/mhoLmx2ZuoHQCqO1noI5MuDS
H90CtpYgDZsxt53OM4rKP25fHXyBMYL4C9MZS/joQNtKGY61NxZmUpLIHhQtHywyrkmFCm822KcK
V01lJIYATgR0eaPrhUoNZN4LD0N/kUxMfDnjneigk+fWEizPa94M1T1QQyFKZNTWnYkwZ2MUzJ2B
BTbGlLPS6Vw0kzJUraQpkXWzsuj5mOLkvaqeBJtzSzAVwq/1qj6GydY76M6w9l/IukzBevBwxc4k
MMkIyU3be5V/CocJFER1laqFkBW0GwOJCNzDfUYzQLrwkk3duq8txOq0eLo1amxBbtXOpj8WWjOx
hk60DpL22fFPA40mm0fGxlSuoGySjBES1GycBcsI23eKwN5eHX0GgRRV1RGQQe8UryRHzygNr+IZ
Rwuo2bB9uIM2D8x4h7MKMG/u67CDdb5rffbwX22kj+TuwO+xn+TpkRRz6/+ihr/HhIJbpZyVQbED
mk/y53Beg3imFX7B0o+bmHiesBj1HTYFLy1hnUIHUIxN6v67zFttliu+eKLtk9yU+r+4QoUArgJT
QxXokmn+ivuC1pZJhReG/2svzt0EZIKjY0Qk36g1e5lR6iJOroSJIG8Q+ZyUGvye7AdX56mC0Oit
9fgWrRCjHPLYhaChNSs09SVT30idepsD1hYGzoUVQVmvWEJcrWoVSezqJQq6ysZ8rQdHJNBG0YTQ
P5VK2E00eIm/fZ4yFBSb8sa9I9Xm93ahjNQA1dz9CLIt0KN+e/XTdHm6osUyb/0XLT+S/mFQcjha
35hy8rMJSmWUdXBIjLsC21L7HgwTM7wYrIqGbZPoPcAd6Q9qKxMHFwytQUUikgFEmchZ3bFndpcg
uIv2V0z3ieEx6kEy5b7fz2ckeQRzRdlNvNMDISPaupYn8QFp4vf31z6KPdBMofNhSu/XBVS6IRKw
N+Fpph3NvdVNQQvCoiB5b2dOqLrugXrrl32Uk1LuGa4W5dAXrBdAtL+64Xcj0NdSke3LJgecn7ym
0wnRhPg0zI8uM3gYHJsQgtZs4QR08eo00xIqZy0YGqzlA/5zUJlteHurG21gm7HZPFrWfazMUPHo
FR9GMc3NbOuqKKlcqPVukSzYz2m77N8DQarzHbQr9UpJpFU++OzHSzrEpBrZEWtrRJtMDRKBtHjr
O4+aO3UYmm6IHI1AYMpnMNNcMykmmjjUzMl2+udXyx7fs+h2gdvXlC55+jnBZLtKKr6+70RyDs1P
D/Y7/6armggDHtM66iHI6uGqk14OjIuJrjMIcI/Z8RhnK42q6BPKuGnUvcnK5y4SCErKhiFOEu3d
cOV6IFzSeVcExyya429hkrwJdQQizuycwaoBwdaEo1vXC/T8q9j3gcgLkwy4zDS4XbHk60tYYWR9
zmKa5iGhtG5CWGtJHf2cQiYYxItllDLJEAzlPLOziJL2cHjZ3gnpRVBuS5X7/AW6x9OGJ+S5Re2n
nwh/f8sqPJBlRY3b+97rW3ub6Cs0MwHAWxDgVAbP4u73/hnbZh4kCDgc2r4VO93R90SoFDn3PLyH
vFiSW3zcMP6nSmUyvVvl7d05uyA/gWDrDITU0iTnnx5JZQMyufc3XKrawkWjr+FcXwDQEWYlZIjt
FZvqcg8+L8JfCyaJac4tvZA+sKiDxHF+55Mp1+ZWdILxrtcm/m/6XSXbSJhemBzWooCC6Rlh6G99
CVcGSPl03V2f3pwTy2H+pdrkwy7tA5wtzemWg7xwvy2wMuXFSNbMr3oPxCEuLIpXp/06UK9SMBly
FCQCfM0d+T1PNLi5NUu4VK+CokyJ0+aFQsbD6u+iOg5XvJQRE+cBbi8ki+H3BG+Z3qP/m06VAy8N
QBfdXWkhUGHJHV0SM/kHbBRjQuUFG+c88QcT4ozKKBc61B0ZqoD6wiP4ja/zmWS00iL70Y88LhaY
2TeraU8K5wXUi/uKV+G8YQsZBcr7VX/yFI0JVXx1rArB6eqFWvDhA4uyKMvEBmPNmoXKM1YkKbYw
5tb53t8AvKm0AokYmiewSdFUOQkZl9BUQFUo21JVxP0VzHC+XxSXZch41s9sGRTGAmEOTOlMBlEY
Z8KY3Xu/XO9sgFHYrQv03Y35gFR1j3He3eZ7VNGGSZenk+ZdfG+QzvyKW+TNo67gWl3oNhYQXPbq
zpG4+1+PUMJySaUbFjmx25N3JI82qaPJUQ6N/QARYfhO013v1oUn6Ud3siNrtwNfQOVtJSVZ2UoA
phOZS09ShAvWVjhE1J4qIi8h7XT3fBae4ZuHAHVVERhKJhTzkHHpRB/V7fYwB1hX0A9YI0LQu3uF
9TIb7HZ/RKUHpSHoBrfk+jTL37vXpi/gLmIujfRfKx5B6bSWvxM66eQU6Cxz28DI8EV7bDDdt9zf
Q9INA7RB2zQdCeY/W3vrR7XPBPkZGMLzL4M/kpIcg4VdIqq5DPPicM2KlyprnCZbR+Q9xLIG6OTM
xsHHIADOsOi8I3vW/4J6v78kvnd8gQcarK2DtJB531APwLi5hfj87+yT3US3ZkQniiswlfnnxj0Z
vC7kESbXMCpnQ6LFZHNk8Y2ZfhIyrd0gwcUAmKAi1KfzjtfjfPR7OlljnIfZ8F/OkCN5KOuJAn35
/qoEQ8p1D826iAPMeNb/NhTFQZ/EBdnoLB6WAZ5EoWsCWalM18ku81yaLWPlh44RoHcDemFKsdVe
/WMLZ3CKn9CH2NHJcsC/hm23TzV9dwuSdvf466fPm7iF8IYugABb60amlmJ+/iwmyxdiuSKI/Djk
4Xg0TPx6EDxYqjtzGRbqHgrpGcL8WYMpy8gwNpQ/w/qi7FP3z05oDMtltssyPkvDTXpw5Zocz1Ae
eH6N7XvYZjZdRhOGzH/I+Smb2ot1VkB8L33DyGxRESheO90RvVRRfS0EF8mOc57/gv/9N7KA3Mke
r36aKyvX5QiVdGVx7cbr9dJdvgzDubho1mbhzawXfxIfynJEF6+vqshYn9gvO0XLigdvspbFptzD
oeY3FVARVwfC/i+58lhrVSOvP1IiNv59S2qvwP8gsu+ukuOQM8+KRvoNvyVhcxSup6gmsM53v0j8
XOfhFlpZs4y7ufVY0WPweWRCasKu8k6ALqhtgWNXxhnD/X5aBLXM3CwUrZbXhoCv7kGcyl7uQj0T
qxpP8897gCnZ+E4/kM4fZKBNtLvB8g4qrfAT3jlNqyAMkvU1hQdttCee0Hb9XPWQVW+Zl6RWcXtT
JXDddjzxpmkuCQDh1yBV3k8GM170DrA/ZZz0JX2lkvxU4yT6ygadOuBr1W7wyjpshoq+TWdx16jq
8cvsSLxghhCoxPRYWyrKVoJl/xt1o+WFdgB9MGFI7itTcMqUvccjwJlC0rdfmdakeE+tkj55D5qF
Ql7iXGB8gCsVYjbfqeMfkOa+NC5zDcnBhUDp9wdIif6i9AaJWi+SN0pk7F2Fls5e3nE6Cg2uM60b
6z4EiKq+9NTADmpRR7Ep7LQXUXafwBdO8lsAo3TIB5n72wdfhwV4LJLuH497GiHoR6g2r88BzFrS
ao6LLblperUAvlRC0fMj3FPZNteXw7SC3dClVrBYg14x/4b6EAq8ljtBoFgw+ZiYN84lcGHLFs1f
Md881Sw6Sce2e77PTau9zK/EA+rERjFi3br4iQd6KS0k+AemmMOIhYAPqZtbBZU/yNkQcvXEickX
z1CZJ/5Uey9saqK5dbkyJuP4a8nq9QBVgV4tBqTnjJ42dw9gTo3xXn2JCF4AmTGUluc4aoypAFvO
OaEG5KgQk6ERCGmJfGlwzOa4GIXI5PouL+i/JhmtNvrrRK1XW5ISfaefqDh7uO1PGIAiSj6d6zJ3
6aI8k+Ic2n7HL0pLGUOp7gtH5qSInXE/9IsPH+JQnlEXjtoajsvLc4MvmWASsMWivWqutIDbjueu
EQAh6w9wIurJ0+nQ6kPh0wClQbBooDTvnQlXFa3ArcLKOJE8yA8DRvZSJ80BWR5GxVUUdwVHSWC8
hbTGsFMFWTwaBrbz4GfaHIbHf1YMvnmN7iO4kxNgDiSMj6v7JqKEz6HVMlujB7z3CZy5Ouw2w6SL
yqssEo515r2/yYEHewNQz6i/s/b2u5ARPbyaYXXeEP0ZVgLT9ZJO+DqmaSmrl68U4XLPLc2Nr4ul
ffgGlcZeAlLJLHgS1VWogbIY1wiK7pkTcMl24bLCaPgnW4BTNrLfFI6gFgKB5IQBssu8mEqhQcxZ
Pw1pNhK18MbPqOFZmd7zzat6RkETjPy/Cx79PCyCkFxPld57NfcmWGoIXIDh8w4hZO3gEdWeSGL+
z2QmAhZrznn5f0Qg/aWb6CqI9iRkS3c+7sIr0Tea3ozB2rVuoKo9SI0BXyb/w9ksc0CfAx57/63I
J837aTjeITtB37ApUBRQob/rkESW4+W3xS5FNL/KGe8MyHxWUJzRaoSLhOLeMI3K5o2czhsX5vA+
cBILxn//NbhB+Pwisp0eHRv3G9y2hMQqKeMvn75j56NcwbPNjkvVH19oLqlyAgXRXonm6NtIeHkN
8PKZB/4uQaLQ+rX9uX0j/uMiiciqVVtDcgipNLrQOEOKWrh6aqmfTLCxjSkzy/CIB9X9YJWUSXC1
nqnIbljkk8b0KWU9n7YhBNfYqekANz/JBKN+PYtGPSY0LqP4YzkaTr00K2XtzZr7zIyvXXEg7zp7
Yy04OggvuwZmSIQ+tDvYwYIgvyiOkqjZZziEDtTxTYpnovrFx0N3MfdeqE9IWGJ/m9JAqP3vSpZQ
M8d1FeDA3K199ai0E+4Lg7UkhoCnmfdN9onOOJLCD7ED3NIKTaFp7wQl+KZso26mv25+nbr468P6
MypT0x3W2fAxJn7MRTxYLyCGd4naVktmJXyHKT+jPMSb4a9ptpF+1CZZq5HRpCayzAgYW433f/hi
+e0+TWIds9BvrJx2AlxhEdpbZDwshoi7waokffciqCF9LfspUkeWSY7m0Rmq8yFpaFkECFdrw9vN
/rFK5JcSJxDPVPAsy9SFTAf4hwAudxUmTiTL26xkeU7NhM05nT4kR2G3Kefe72DjBMTXFJPWKLpy
fnxZQoF+trxLt4meAE8eblpEXCIVC4ed5NhQArmJ6Dt9KHHDBLstF0v3bS4EyIwjiXakotaCbktM
1LKn8AKCn6QZEfvgcPVDbC7jtJPaApwysqg/qXhbMjWu+JM4mryFI2eMT7CketeDC2Sb35z0EZ2g
e0y+yCLeLRV6k0pq2AJp2dLn8xR//ofXJoNL8wU2wOiPld/Z2dswjjZQzag+LvcrOfr4Lk6L1qxr
4unhTcvKv/eHoM339cTaE04YjHDf2JGUM7dSJbiHsWFM6ZsodJcR0T+1JwdLRzPgahkcu9BEMo9a
cW6y+zzu6f1St6Drghq9W6HWikmpv2Rw9DT4hx6JsBv0T5kgwthEyO6J7X2xwR7UbgGjPrzUtazU
wdAWqhl2NVQn36dj1mZIamUno5KbUy5KbDohQFot9kbBLBxR1MLrFc5QbvrxHUZhMHlikEegnALW
mv3Pzdq3A6iHhxKQwGig4I6HC5wTvLij3QAa1lLmIOu7eV0ymYkQq5lY2R0fA0wKT3StqjuWc27F
UIeAGd9WPyoXzf0FYIBvPd2Z3lWxv6NdqPJ8wlOWXnDhMZ+ilMW2S6g2M0i+cIzDyOQUotW0i3GH
4e0Hr+G3+P1McCyLqYFAnao58bLIK83yOpEYiWJVWsrd6zMlPh+jjHnz5T51mE2ZqkZ/pUOqh5f+
Bu0lCVORJ3HCfxiZypOu7TTVS2ddTlf+BZh9xauxkK9W4XFMZJ9iIBQvz69Pw99IkWqALM96Nw7a
eDQ3Be+hwt5DUG1XxdDMEhjanMXb9FBFFBZ7yKXN4tKKTXl+s+dvrD4MMqvEf9oGhal0RbmyYCwg
gODyBd5mFDoPsQMHBYrzJ4rRhZC+EqpC7meEfhKk8IlmJkWNODaA7RY/VQk30YbbEJe/XRXzcZna
j2LuJ8eN2OTYWPASD77oN57w/s16usdk/llPu3SlZDfcfAsP73xEwTdNDYnNrUN4pwIEit48LU89
eCngy3J5eqTwceSWRPKGMIqA8dRUDMFHnLHyg7fdFEKB/C3fsbuS0UW0D5OBOTdCepjFGTmTButu
yMWX/NZf28qDwVgkiE7Qfzu1o+sRdLFP2IqZ8h5qEOPKiW3mLL0G0TfTk7NOrFoXs7OTTIYUkj/P
lFYhxtRDS60CINJ8GdpWzAEK6aLiFtCOsZud0AHCefcmvQXcWFMZsqCZx3NwNTMnI/JCO9qk7vyM
+d+XNxsgD8dmxWGdvJTpoJQmV48o1iNpV8qMjRrD6vrNFeSN9+W8ov2QwWu3GHrOQpPuQn1ZjD6I
EbW8TkVAVYE3GQlNYksKaBjh3Z3VzNpGMpnsb0D5KrmED3uprtAqnU1wx7iSSdjtxbXY9B3JX5hc
ompjujX4DftaobXJ8c5QopzBnofQ+QuABEA/3ShuvPd86tSakVkindrV8akd53sxmok1NT2QRJjW
ESqRTSpDODVSqp5FHs29BvMaiSHr8Lbh3HiMnmg6MOhEr8Mj5xB5/OYk0/5XjJvdVCCBNCjpw+Zm
B0vsdjMQs2m9tzoBnDwMIxBn0cblui94aSr6yLvrGaz14wYRmaFDKts2HpQrB+Daj5xS8B8CSsNC
xVXVysQXAoiCnUkIDUoGKqZKur0I1XugPQxMh1LwN5Ad3wXQsqawgjHmTFvfgNwGv/mNaqd2Nmr0
m4Yl1522SVGbn25jdCgYHLknmEUtJ3IOdCFN5Efw73vJeI7KEjjWk/g7zu0v0TibJBjqlSdsuY8X
HDxWU+9Wn5kErF8MPRigJ97at+OqsCedU+DYyfz1+DzDEQwVdrWe9qYc9RADlonlEeky9ayEup2p
M7Z2cHaqfHR2+a0zMuVL1crUAyQURUptm87502FsBRGWrZBdnGCH5kqM/yCckkIJWfgubETBj6pq
b7s0AJsWIugXXBLYDm+scH1XdYnCyCRuPWLzNWcMJnyFV/jupGdxyKUCnO6YDBmUZd5AhtZ9dC/d
vPnTtBeURDurbBZY/5DOEMReK9cx6Gc7y96tQQotlcjwM5rIBNjWWRGhX8O3Ym6qZF6eofwxi79X
X96LOjN8Ogw7uYRhqxSDlNsr4oXsiHgNG0pNLJXX8IlQ2+uCU6pBFfADxsL8ifmP72NRDGyFha/r
XHmG563gprNbar+pJrVROL2jk3W4C5wn/S5XHLPwzpC2kDmkEM7DfT+DPVHvwxwT3Ix60NfGF7Gd
bo4i7lvJgHuYnMG4Gfu5fei50WzqE7v5//aZoLIZKYHTpl33iQzyKWS8g31BTiizr6kAxSArS/VN
2EhWQERK4qfebfO3LkWxmmaT9rW/BQ7uJ6IPuhRUzXQaI4I7gvLDTDokT+Eje0OJ0TbjSfEh/5JM
KNJgOmH77qEdiLDZ9gXKuREIU+iksDo+PmnboIqFFPH9+cbYPEos2RjnLSm9KYrTthK2xFk9N45t
QfQZpIHABvFLQuv9qKA+SYy+/+x+ubMks+0VJ55tD3ee5f3qjZs0zRQr8+t7Ajg1IzD6p2N4WCtc
g7DFonCGuUsbyF7+onYM4Hp2JFRukK1BaQyMOwooQDjwaYC2bZw+H9i//TM73hgiT23vJzzTUa6r
nQKpHxQTt2voYG8DzkZ8+iCZzR411pMXUM4jQwsbSud/WJMQvV+dxSi/9r/SKUy9g8pULouzy6Ts
y+qktMAO6+nUsEDyYnW5K5Cxc63XlZ2/2njZxukcDfF+hE61gap8nsg3m3x3iPPrR7FmMDDvzd85
UhkLcEIZYJm6hS+TBWFn2JFzca10nfGCCMfv6RWW+VL9oQIXwmPZgWPsVeGGF9PV+dx7fVt5iFIw
Tr3ziQuEqQ4by2u5HBxqx8uAbB1yQWyoytYnY4LK5WtuZO9voqqnZt2bqT94sEhg1tqlgDaFPb2I
s6UFLPm7UQAbreOz2IE9txCIzXq/0UU0B1Bcfnj7cEKlTQBGBJz4fPeiy7SZtQqE+u3n6Kzv05OR
WkDDT+4UMKIvfPBlimRi7n7Uvlu6XGCaWE96gxW9gLSY+0u0f0F/Fnep6IeEwHe5WXzzNZf9rNzK
m+qx70Gxdf4nPvmn6F+gkw8xPLEZVWFBQjllJinItZNruJ19Hj1Y8zKi4V2slt/k7ztaKoqf/FeS
wTDVHPsHKloQoNQRkU5uSn4Si0NN2JVQA1pe24RSA9T9yTG/8FlEJ7qdCbg32dbvVQG8mFhVKB47
IN+g1v4Mr7QomUAYxbNT2HkdPBaxmyXD+IN9t+zOlVuH8HV9NzcGbM9Cfw55nPEAOaEPlcMAXGZ5
NlHUt+rb2k3065kkKKbFZRTlGwubiOm9ZQNW8QGK2UNE+5cDdcnNAIzW+ZhfGwBS7bWmjTrJzG/m
8K8KILs0WRqTmGMS489Wg47oz6nCOQHxSa1O31D6rob0jeAHpfs/YMLB4+Dl5puD9T/RV4mRzGqG
BzuwqXrqNo/glabBjvezhS9NhPrFdBU6gX8VCeh0XxEtFlzlSHBl7p37V/+8Vh7t6M38Vwa4KdPM
KifxblUs6pmSOVerFviLPMRohfEhcRVnquj8zZu03mTExA/qskuqxurXbBFuzmIYKFrdmMiJnNzA
ZYv5B3ZiLhLUhMfy0x2HCF0h0i1FfnNvrZy7iOsAb+NaJ9xWAc6MxWIR9zVTUXHbFMBVfTAnXyCA
2uVfDUtdgoyxaRPfi0qiSif/tTwY4Pyqnk7li4BK8y9MuziVYZTa1Cq/z7KLA3OOzmOvu/91jWAQ
TXTOZOGDIiGvE2hynOJwlLa8N89i+wZxpYY+7sJPPgeQRhNY5dW1TbBK5/hhcapIhG1sSTKtl3BQ
SSaQ+S9hwkDjgOCw9Xj0qd3eeK37u3g97H7SXttnte3zNSfhYoAfs3AT/+BOgGKNzYmA4xZyPI/M
Zf2LBtj+tDC+oL/Cf6VVRxlS/EcGdUE4sweEfDjWUYgZOZBXNzshl0mUXoGhupdZl6BXnH2oMyc6
NX2LUCqSDe2CP+FuuEV7daxq+JIClPYq+BdIpkIETpuUCNEXUVDHOIB8eAj0BXq2DETWT/sFnojK
ITmSyB7ARioDxcXxAPTw4gdgthZuAiDurW+n+moub7300tyztdK4Y2p8WKHT85Q5Qq2qMA2M+8h4
O9H+Dx3l+ICqvfdQegdAWqyyB2inazZOibrZhxz7FrQ4Y90HmKk1k29ndWLHF0jfb4IWcTFvXwQA
/OHdfp9OIGkxqmUjHWSjrEuv8JmHCP/mBvWZRhp4NLn8/tv6GLiB3X34w2kggsMX7iPCVYbETPm7
LUhTyORb7eCrou0AXwPR2nDDKpUBlfnkjzN4sU7mZmKTzE/avQU5WLGSVkBZfvFigtM6TnDL/s8/
VsL71xyVmBTWsKbdjrnGtcWFDWAL0Gf871ewI/WYOodo32GBGgnGoATPC36N3S5B6fHWixFLFpHu
DJ4uwuDC5GIjP2lBzlbQsvYsghSVWk113iIIjQS9rPzaHn4fO3Uh9dazLXNqI+VOt6KUnpSrWql0
7L1BKu9exq532Ao7TULo5Al5qeaEn7GToTm6/LcrZUbRrCPRmEO0QHZ8BqfbMR3z/IME913/M24I
LYiDmyMlPMG3ebIgMkvk1m+fYVUiLNLurngSNezSE0DouEEbcwSQgjBG02shKX4f90fRYlp1I8bD
OScY+IlBYzjXBLffLUaax8O4PcGJ2Mn66UIMY2MSc+oj2II6OZJtr63TpiK44FYia+B77aNBjCFc
otIsyNxapeXEg0XBXbZnT1W1uehX5RITzxR02RR5/IZoc9giFRWA0rDDPeNcB/hokysPMEHYQQ1N
RAHVcfV6Inmxx25mS0G73g5TRVKbxJ4T5plzLJUTQLRqgj9BgducOLbfDZm+Q9ssjZlRe/MkCsH2
2KX83OfkAX0DqqDbGTmGzTzp7VR18Xq+G+hPNQ7zRICYfTjbl1RGYUfp9aHrF5Q1c8E8oMi4hjwt
CQbXMjN3tUUGgWaQSw/25I+K6T+xuuQbRTa27IY2WrWUW1JgCNQEmspDnBfvLeCHk/RUO0DPz+S0
IjRgDa38sm1F4bMOrWGepJKiQWA6c61C7JGMqAwcABFEJkbw072yLfp8aVw3MGnVONL78szobtoY
hy/XJrVSuGcQzbjvds57XgW8ZkW3q/8AbwlAj+GOHEt1CBSPzxWLtyis6u9W4Gn+wsk0lhR9parG
pJUTLyx+E9dg4g==
`pragma protect end_protected

