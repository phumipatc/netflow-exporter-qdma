`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ueRfDnJVTVCgjsf9cW/beLZdXgzbV2W8PYhczBdVSmZbeVtLSjd7JtPSqxIXv/MtVlUQmj8O5wiQ
UCgMRCbxcJkE6/7TzlxEM21bIye/RqJqYvmBuegIEjX4ZIitGBDUpzqitfXsgB4PANwqMidRUUXA
7+C7d5zY2zNQRD2jZer7MMwCqFLBKVN0ddLirwmQivs70uph9Ur2B1sUy88PQWqPPQIJCFSjETlG
+5sRak0Gty6NT/thkVXbUzjbFDYz16DWJkJ3BhXb86V0oOaI8/G2HE/aWY2OZ3A1gVX2fI4sEdsf
b8CyJDD+OrHEWft89SoRrXyW4N6dGFBUxTM0yw==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
Y6lo9bvHZNAst8AJFBqlO+U1UCG2hpiJnANyYLMw5QsLSd1FWNqiqywYopVyyeqK9DwtIGROXjA4
9PqoiNAua911VH/+7q0cE5lg6Bm1V2JijkeM3TftBVWBk6XmxAUmx1yI3mOJZsnOdsezpAD+/kIx
mDwA7p1hskQJV5KLqcl9EdxOGcwohfOcn5SbnfvyQRZGa/bS++w+QDhzqr8qmbLCuQKN4OQHFIi8
xNF4EQaaSyKDRTovMc84tUZL1fHMZ5tsCr4DaIfeISk8uQY//5CgKnL1X2LFu+LhIf1S8CbLUCcA
zS9SbwhoD56GpcHb0vE0gYdboqYZyMDlBP+TQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
ANRA2pgnChCFrC4GCt8TmIAR3WF5eNXiSlPFUoyr0EnwkG+i2CSP9Ex2yxCA9zCzvUyYzW4UzWoa
6eAX2jJ5aA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XrtMaZmHIO1eJ1MdQhRiFyf8jEGXcVlCnXcGA3XOW7d+M3R96Qy7w8SRMm0pY8KBNehxBP/QY3mi
L45+ATjgB8bZE4gqm69H7BCzaplHL2etTsDZ0ySz5OfWRCb5LXhvMWNZeKhCBs2ZaH8MpdRxYbb/
8oBaZrTl6xExshAfmZmLsTDmR4j61QPskp1UKsGNrTTjEzWZhzxIdXHQTaS/l6LzA5LQRVf/+63S
vVz7yzqBkvTEm6yVSnZi/goSgr5RWT3Ap018r7YrKi6kTznVLpqmjR29b9PguXZEicvzek4SugAQ
D3b3mv6pra3ifGJOvWttAUhwXL2mWQ7TydR5lg==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MNsNKTnAY3yNmj7+GIohavN9Nvz0czGijXQrfdyNCZE5ACsLmC70nFVn4cWE6o1r2m83Bx5LfXSe
NV1sqHaepJ/kl9RvryoEr+sB5cphXZ0i6e88d+VMeS9uB8AJ2/jA8M8crvGcvYtrr/JQ/BMF1xmB
1WJt6iL0b2Xupd3+XwL5ERO1Arr6Krod3z4xs5GS8XmjyiC/Hn038Km7TTn2bsJ6zHcYjjpGk00N
gfwLsWw2ph1dgUF3pByKqFGBVo9cWeZCkDoRYZ2SSpAfXyIkT+ujjZyNR/USx6Z2uj5EB5pPKG+P
UOMErgqBGRbksbLGzX2LeH8bUUkcXULxmdJyEw==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
uSnQzEgxVJxTIOMuFtEbKG7pOilY1x/3KNOOAmQ6UgmMlK+tLKd2cM3UkuLdtBmheWmqq06+73QF
ryGJMIz7EzikZ7zxKgNfDJlMuj311U3l3cuXI0gPH8/QBgUkIntu0uPE3YQ4Ez+zcscRxcY3bRrT
Xv/9vs3xug87DKd/4Ws=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
p6U1k7BrHojYcUw9NFu2p/ezzhPjBXr5wzsvlyHK2NFlLjukE6RxuHdUFVqESr+6ztO4bkYjco74
7/a2yrpq/DpY8lMd01C5mDjeccyWG+b5tBgv0p/tLV7JEpUnX1kGE4a01DTg47nuFn/z6pIH+8uv
rkH3TSkGOuBxyOY1lskAyroKGYjJvGVcQUQoY9KRD0G8HAuCyvsWv9XuUk77oNacq64wXgvK/Zfb
GT1PhWq+e3tWwAE2UbuYnrd2n8wm8d8bdaG8k3GiagG1n7K9pumvumkLpihWlNtPIw+WuIvHkrTw
r+qSAG5NiRnbC/dRKTLqXBWrzEBhkkEgs5rXPg==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A0EPyLdoEV3wJ12CVlUhW3GAcfnXV0eOTel/mZgyw9cM8WONWaoekBimgcAF8lmdNkcUg7+V5I6M
Fg18gqYorNG2daZnA+d14SxJZGijIpsOoYvPsJbJS7f/IRKDtoxJNVM2HlK8qXjOe9F3Qbv3JKwW
nM2bCpV3LZMUbxxEfdXR8W1N9+pLMjYadXiGwaPvLyvvSKwAXr5YLuJSebi9fawgGqGHNdGnR/BM
3jZXrIYWrwfHS2EtffC2dBiSJXfnfya3bxzA5P2wHYfBjUbe4jKjR7wVivXUhoM7j/HZlOoTsTbh
fCtuFcHwiokcNwEpZ5t3slqJNUMVJkV1Iq2Mzw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ERppbtnCDsDi/lI/FMSfBZZcLkFJP6R/h93nWvd+m8+42TBCKidNGYkECNbPfOOzefMhBlY3MxZW
UwoAJPxq7w8iI3sarVZ4GkfP/DwYAlo6n22WIAQuymw54gLwWt8pnmHAotObJFU8rhAvq12iVE7J
W7ExxKCa9uTWRyvwbfc=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
fSDXJCEk67Bcq6isp5qeXrYlzjgu4+pFETBJGt1yRH+rFj/r1LJaWQ+FtufDJXAzTDPqwzxLkVel
rmaix6wRpkJOgH9ykW8YtYVsOzyKnvLQU0FhbDwzyjskr50UsOjSQCyPoiAFZOw2hOWiQ4Ws0YLD
Ac4X3WwJBOxDuyJ8V/jOYD+A3/LTfDd1e/4Y1QhbtLxN0yq6VLqFhNApOfmW4bqY+Dum58jzIiw0
gnDcr0GsITgOcve7fhsl9FhvKzLVJFR5g7iN6GzoRiAcw0QPpmynMoxJ7DaXrRZE8bqxVgTZ+Syh
MhEn89QbJyU13WLPkJd89IuY/XSHTrdYbLtOhQ==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40256)
`pragma protect data_block
T2Cc4DuJKhw+qjqZrv3gokLllpKHh/LsTCFQG3iixDBV7zye6auZ+RtpHsL5VzuBIbu6aN1nrHCs
c8MbggTD3qOPSPQtKkpVsqoSUyQx0Tg0wnuNX7qodk1y55ZJqZoDPVxBGXlD2wbFjc1xUjMidkq+
C4BCLcUivvisjk1nOgD7jzR5P56LAp750GV34i3YtNOEKtPcmzaAcMBiHH4nrfTP4jPTH/8nbd0I
BwopXf/0K1f1iklr8ol9Zslx4NbkwMl6G5C+ie8K6E87jdIuil1ly46SD68RiNXSTIHYtJ3hfv7v
hpWVjbAf7YwAIEjUX4nB9vg6E+xaYhqlX7jVg//Rf5PiQNvYCYlDiktfwz40Z8W7p4Qavsux01Pk
3rlgfJVV+csYHxWhE68zHTWH3BYDLj6fjon02vFKQ45daiIkpy9w7xWxVRECS7Eikwugl0OabpzF
Y47Q9jOyWPzF5g5kgf8YMnQyQd07bIHVjTkvHzm0LfOPODAvqXmfDtSrhr6KcqnWvu+QFjDnAo+E
y4L/HIqWcPg+38SAgK5b20caAnGbWjTx/S2FLWSa1SEnGxFuF3Yng/IX5HAINKvK4uJrlu+c8TEn
1AFiKAoJYwK2tkjKAlmjID2e62mmg1T/2X64mqcbTukgCcdRmfE9LJpv/dbAIV/9MV1zPGCtGy4S
ilr4wL1lJk14J1u7YkiKEqMv0gsCkYwi9QBFg6iBvIHmIIhR4VVLgbTqg3TZfnyEWCTwcC90xEbf
2IUxlYQXV0swgMT2oRE0MbcnWA8cLy5mGFus8c51/fch04juU+Dde1cWNVXtFB9pF+th47gQkcnb
ydBg3UXEL5/rj24ihkTfuEIXaMEU8SU5jqZzX6z1VpYSzbht2J7XaLHlPBVxKLZ1OpmBZs9KgL9N
L8OtvUjRSF4GJ7mZHsnfVIJ/GRKLONos/yijVi8PDHhZlMg83Hp5YhvhS+wBCpoCadPWd9G002eW
4ffizHkCZZh5YS/pRn/sBZdcFNz88q+yem64vQI901hKq6HgUa/SqkH+We0ZA2AMzD1fswUnSu2Z
In4y7/bF6VC/N+f4MOJh7M5nSAXh5XOyfwMR4hepvKAoL2pTuwbGEZ6OVq8nGQiOHYy0a4GKVQOg
C1TFwNULJgrc2OVkUxK+13cv8stAkE+iKyXSTFAfBlO7EBScKFQwVPA+kE6S+r6CBehpAmKGjsyE
6l+1swLN2t5oI7D475Jqn6W2w0AvuFE6lRYrcOZJy1k7t4Cy4YZzLXMJ6w1p74nNiSqpgWV2dEL4
rMQd0Q8F91DJS/X1TaVt8dlzOEFoSiFUFewE61/XTipNYkv6V8X3ZUbPN6Eul2WvhSvVsA4zb1oV
w4Tzd5Twa0ZPD4+QQoa/UMX6/7jGUO8ezvdDUc0RXrD4mMBSMFt9N6UoiPlTrNjC4gLILpSSbJk9
IPBTCDigvvbc3WMKjFAgriJ8Ky/g5Fe0/rr0kSHVtgwnCTBt2tFqWecDxkH1sVWohDqvjOU3KCIj
LMPUaykVV9wpLxV/baHgPVicjtn/QSu/dQg6n3VG7uDsUnE/zDKQ+FF5hgKh2A5md8Qrkzn3NaFE
1iVFtrFyAaaizZWKQwU/YsDqj/qxtS0ffguldsjquMQCyhLFDRcwCyWeyTSu5sdnIznS1ooHcf51
go31AVqaFrLYo6SmKabufiDt6nI9A/BKpIctcr/zpogI1z7G862aknlNKBcrvxPhzy/wI5Vi6LAp
3yRXcZkaXV5vJ0EJ4GkY/ecr42KwCnKdPEaXChlZ9jWMDTtVhkKg4vHmyCEIzHfaF2WMNZ7QV6Tp
9eh16TeaAubird5VqP1nEJxnl5AV2LXSnX7OmzFj/1N5nKyGSYdcT61CB0QC7FS2StEZYz87roBx
dJXJojIV0fhk+Ik7qbPiT8Sgc0Espx5iBwCh8SyLDmLfz7/Mt4QuuHnmbvDEQ01KwbtPuVhq2CU8
63crcd4c14SceMTg93f0wruuYsA+fciaxtOgfdXdPxjnZBYFCz/IP+gG6N/DIZFEEhk2pBxi5cHE
nT558DVnoSthN6UYFWJnk2wHGE2S8PH6FUo/aZNddTMzLm64qaYbHEvgiV+3Q3o1qol6GcxOKNf5
Gv3uk5lUJKWkpvBReFQictGhmbcMTstGQHV55LRDWb3S6XCggxwpt4+50HlGvCgfQqS7NvcWzLB+
APzQjmjqFpiDlTd1tqT4p2YW+zGh2o0z30ulHNuW6c1uz2DAXUosImXcMeZFk8zESzBXLGfjsetu
S+XFDmD3IyM3cDMi3wGc/yb2VF5nSvuLzM58Qy9jeF4ygrFyvoRzmxHHKBO5Uum2lgQ7U6tHzKPh
8js9I6AD8o7I8nyRdGqCi2VCAfuRgU3GnGP1uv3kr+Bt+IexogIEynmku96yTdr+tTeKtN9EDn7r
KUTB7TFW9DPC9ncv/y2sALjj87f7Z8pC3cOxLH8XiTckxSiqo3XGrb5ljq5JxkEVtXCowndmOI3Q
IWHcr9QlrygZlJ0B18pz8XOUA3pGfhRMK+6RoPI2iZNFx6pE9k9umtqim7m5l31Rk6B6vIhQfD38
VzTM1wI5YM9S3CAkfrfRDxUCk7wvlCEajrYR8OpUoMlYTgRt95iHr37/aZEuJWFm1K2XiNHXFLmC
DvbNkbrTuS6+2Ovi5EkXy/YrtcSsYKhyAcM2OqDU+hlYxUpdf1OCwFSWzQ3uzzkdyQjj1Ok7i8VV
hI4VlJzObvR0Bi34wvTWnxKcX0WY4Z/fD7Y+zUfkCHERQI7mB/z//ZLd4g2b7FUtA04t/DDc2LaZ
du3FCFYffValCFwzo7raR+T+o/LLJgSH3WoEEyfPFony97qqnJqqPla27JfCLTOQsRv5ZsiRtb17
JfBg09MvoYzOOh8hC6+qTKXyVZyT+MlMaSgMxtp+lz31dFhNc7YbrHeHcg7Zs15ZTifoTmYoywKa
k9pQdW7bdAvb+IRWJtlIzZSRSEnMUyLjMUaLmejkW6NMq3JhfSD3UDw9SrwslC+Xpd4ca0o869yk
4Ezcvgzz5aE1yjX5bXGT1D/tXuzl7QB6G+nwWCVlhkco88M6uKrP9c8P9tyLZT8MeBbPvD/xKnc4
DXKoU7Lb3/mGtPO+9uiA7mqDIi2t94W3qmE7rf0iRgr/pvRHZYCfTl2kUhj+8eA1JDyNZHbMkz9P
VJUSy91+ZpoIbtMF9RsLvxuNjdvgsH7F057WGx+aYTyRPT27U6pZ+4/N5IY/tioeGIEcZKAQqwkb
BUoQoUA2qDs1+MLLVezIS2Wj4Kg2Z58yq3RnFJrDPoKW6gn7Awy4uJFMZXhRl34Memb7RfCbHd0U
Woiol/NsdYaya+erjPKbI7tySZpS4uWNs2lVFazJO7AFPqRDhx8qLzF6D2YLNfXkBkJW+NNAJvF9
YJtXZjxZA9Y+Au8jqbNDt8ym4+jHJWEBIYzGpPPKne4fJRV1XpeYyVe2DLbDPz25nNa5UMpLzckg
G74YD4jbMmx89KhqPQH7jFVpAJQ87qchuLNlfSHDlV8MB101mwUMvjIgSp6K6oYEKtCoZidoE79/
C5/2nyKZOqYGvUlVvDWvGTYHyMXjufH0TVHeSvrRKN1cVHww0qGGFaxJvZHMXUeGt+cwVirIWK4P
c8RF5QNFxSKp2gilN1xfdlLgPLGGXj6Q7IcG8lTgoEbWo9YA8QpXC5VH8m0jwXbmVAtVgzyAqLc1
dDIGwVa+T1jKZjWisropRvmrvGVSGQELqhm1ZIdlXrd/WaddTOtpOmlpooUhChYogY7XYL1X0R2c
bRzQ2j5BdPmbpX/UVTMDKH+t/n/no51KN8DkOC5MSefJeRMyqM1Qnf7Zhdfqo+7uWSL0gUe56mpM
fcBp+fiqVb1QA6kYUm9MmpdF3vlyuT8eoUuIQ5jiGsut0AHZWyVoNnEPGLkDBlXFFbdohL9sWxd8
lmf9czHVyZ8XdzF3Gvk/msQvOVweJRN/stIiLt/+Qm/H/KTeNAjCvMMfy8t9W3l01Bb7G/cJNXzv
xFSv9cu1ngX0EP6Ta/kNP2e+UlFo6wKrtlFhts+oI9kE+k9g73nCx7HzmZQZ6tC2lqeSOCYVA+VO
4psh8dOkF/Jx7qrd4d7sSRJATuolYC0ahJ8JVDVYxnGirMlNjuRVeXGBb9H8edhIdD9E7xjbA9Tv
IXVgSY8xy86yZUnhIYeyKnZryhsSnsRD4Gg5LqkGsIYOZROtHeb/cPgsH6Pwp8CkV907+LajFvXL
01egeAl0mik8UkgrjEtyPMcDhuqJHuDUjgFS+Z8p22vUkP8xeqKJzDANT38bCAkViG0IKm5ZgOh3
RO3pKuSiC0zEz6bFBzyhSzvB7l8el5GyG3O7Jre7LbXjdQ0epBj0OJocJGPQiP0V3PW5UWPmcQTW
uatnPOZxuwsc1dtVX0pDscfeWQmLiQG7MtCY3FP+4Uu8E2iRKm6Ko2umc5RFXBGiYY9icjn4hk1U
gY1098+qzfOLL0wG8ih9EKhrzopYdpEJ1rZiJZrq4ucPQLHaOmYmKd6PH8DCnAgkkLxh+NNwX7pt
yVZnvZV91AkyH+I5iZbK7OWW+UoToJgjBZ3xM58054pnlco9wvCjbLoYY3KLG2O8aFfVL2ZA50Bz
CmCZMqg546gIUyOYFygKhGV9dmVg9iGt/0/a+CvnONgjPHVvcmsOVLMEO1E7kKzpmpMjkboJAyQl
11YuP+Wo5IqgpZfQ91jjy0CBysFBZRdlTgUH+VFH22WaHK9JbgGGlS/hrGls2OvL4c6IFMmGqHFD
VwnzBGgQrrwuy0AmZGMKa09kDcm0CMjpMYKUEvxwcr0lQCfq/hLtERb7aCy4TM5OTRXaPu6C6qCI
SrCQvPzw0xbGZUIN3J7bMN+ALTQ5sMkyjJZ8klcyh4h9T+D7bhJ8MvM7L/fAvjnWMCwl6PyWEWaT
ic01WPj9g6n53UPiCopQyYXeEMURvxQzi2NTOtYZl+eSz5Ib9hy8yJNnWkRTzk5DbwJ9O+j3kh+t
YkewLI4vjYF4/0qrAGJhwbMR+0y0wqnw1GNrE2s/8rfvsKSncS2iFh/20EAMtbpxezacAEsmKJRF
nsVb8z0VHDBpK1PqJpi2+TdXL7iC5X8/LmCL4KLa3obWsy8+NDbywQQqZYxJMsE9z0jBqODNPg+B
nMno2wn9MliS+pbqaQTVxGq4Adygc9EOGssqRPREGB25C712ce+fEsT4qdRQeoOeavECZs5YFruN
yZSrNUkctTDHt/SSJXbxHPRIPHiuxu/X+kgfd9xUYx0KAYBLOyH73juEjQwLJBFDBkJ2U+LYpUR7
wT51fRZYUL50WMe9f2rUYVBcjy50OBZ/bX1joIFz6PpiXyp5IztaZMvEDFb5DvO2r0CSuhLc6Yp/
1hQo9dqJy1+3A8KYqHgYREM9d9lh6fCFVGizccn/4j1hkglgLQwL9X75kAqobwSQMWARu5ED0sK5
HxQFAtVg9BsmdWV2Zx7LuWtug/K/V+i/Ek2sJRuj0geIJ3tDivqZdtuxZDfS4ehJg56Q+HjWjzkV
YRrukVDrsCjmxZXo83qvvGSaRv3AB8TkyWBaw63Wh8Kn6OVf+OP/+Af/ohkXD8yi/yju+++bntlK
pcoVN7rskUmOcUcrdDkcNtIeVdMypEpIPx/La17GWp9cYFvql2RoOeHdNWkH+58dAPVeU2HZoryR
nJ9ZCdB4amN6c8PpI2KHVZK8X9TVRFoYo/G4TT1qhlTuvS2nqasAIoarSM9JG49Gzf1sTWaSGsho
Wf2QXd/7R7XZ2ZN9Hhq4AXJTaskEt+V1wnn7qtjKhDLm+fNGBrTF6BClgCus8HBXMTc6HvT4KhZz
L5joUEfAUBWnR7vlqEhDorTb91RE5MScdAL7v1e3WilSw0RPkhovKKows2twJwe8yGKM/SVdALMF
EdGI1in/WZoTRiGPVM37j6ZJIXve1N2CEuSUv7EbF4t6FynKXqI982/wOTwKIkK1z0Zh9aMjeTxy
iC5bHzv/LqbYYLZV1e4IUlEGXacQ/4sayHWgh1vkq2BYub4nRf4rdWg4mrh+BOY29ikLeMTrB52g
eB4e1iiJCaV+HfgjN31RJzsmY3ovLEBlsTGdrpWEtO0UbGtT0bNHEAZF3aflnnA9VGQ99wM4q2UI
quthd4rGbfq/sVdCrpiuVD+qICqHy2iq/fw0xjO+Ce6s3FXMfSeNQ6MwQ3zrnNGCcmmcx05A6b49
eyFFDqe+JRkdqcKqGlpSjfaLPoZIWOJDr0sYsMNSvqGPcOrnauHL+buHpD1xw7LU3btz126/lx9H
TGANB9Mfi22T7CrBMnbJUJ4Gx83R14JhRidvFmxdZYQEFp+bny25QNTxoPl2ZojntVK/KaCa15jV
HXI/VTamRz3DtoN/iVMw+kEPfA5PBgvZgx9v7M6LF/Qt2Q/z6sscj7q8JFSC/1wcAKVOL0WcsuxX
uSeVdpS2jqbqbId/NYXowreA53vqof1GDZcub0qRXsztvTxnfBhn40V7uls5orU+sWNVUaTGprrw
58pmXjOoVOpbWuUOcLkJlDkU4EfRGevWri6rY+vF7w9LPR/RArkfW8X7rXxD5VmbctxbH+huDFJC
S9Dlwgm7dHpfp8T9IKzNL/d3ZZLa3J2/dFlTP42lhj8zvrXzjJBSEV2vnNalU8l3XByqY8Vj56gZ
/lAyTyoLMLlVtK0nvBVe0/R5d/T8YHEk7WzjLCGkDOPhB2h1bLMFWJv1IChjcJrx3wK32K1JLUxE
sORYo0MndLZwo1Wg3FVyugWAjxqtt3Fl0TWP78J+lsUZzweTltbHGECpfxrPWkPuK2nE3TzuxjwK
opw+DraUyShZDKArh3x5tguzP1eX8d5GsxWiY68lpbI9Dtk3mGIoOLL1rOdGvDJb5wzK31Y/MS3I
e3BGHpwRkxrFdwGUL8F7vu4KSO2E972OlORcbaSQD3oEtFC207DyuQIaCKf12s/iFSV0tE26zvVY
jvk1sxCp//bA6gq8ZPMcyQ5FL1v5L3DS5tG+TVwxdoxpnjUCR8Lxwz1HUCHRFfJcwFY5l1+FbjW/
oydB/q5rFciGrQMaaw8UZOGWwaqiavWLswvx3uF1Rh+2fqiLyfMQuE7mL+8i647BreGWbiSGwRox
zwy+p0Vp2VQUHcFlxIOf1nP/AgI7fAxEVLbtoCKo7bsZ6X2bUsmJ91AUtwLSBSSneEdy/HMLSqTv
KhnJ9+Aovb6vPSxlscpMGu2+nR9HlE8Mwbv4/k9S3NXt3xuC5FfjgJHs3/xiRgAR8qSpDsNOL2HV
DcPUIg6fpK7BNsEtlolCEfVFjwRgoGrBucPPxzoaXcHvi0C2YKTANoy9Gff4Oi6HguFdNAuCYY3N
WXpk2+HWPV+Lkvg7+cP6roj+vcCFNMKTMaHOm+yIsqSlj9IBlcFv7AEyrmDvxIMCnwwvrQpxOiPw
mzbuqlp97lCUs5opIrj3zyteMrPT0DarfRqEukOpaOhCVUQ04jYIbqvGyu3FWh15lTOhRXPXyq54
foC1KfdNxW8gp3TepHE+KpzsARzfITY8GiTB9loeZL06W4ak3aj68s5zt/7t0vrq2LxGmqkYy5EX
6JQD6PY2hWjE5tNdBSWJUDt0Bqj7iGaLvNiWz3GUbqxX1aQkv/bCWXJVajauR8W/96+4oS8Mg95U
Wdt5ymA1vrX9+kMQFPDkglhh+Ym+xk8cX+WQmZJAvwITOkQirtMkx9PADc5o+CEKHrdDSHakOQlT
/iyZQAKRadCkH0OUlIHl32y8SlSvXyTXJahIte1g38JY0k+TGU2V+fNQh5CLDZZaP2EDk/nMDl0z
fNp5Yq+dRK+wv+l3p/dQDQkCj5StKOUXLBKuyDfolaaep3MmvaB0tDa8aZ8j2XBja5Z2TuE6tTCK
lo43uCMB42P0s/dnG9LZWGYxJ70BBcNhayU8glvVusLA6XxsZnANPTVr9Ol9WUm9cCPpVEMM3hBP
enVGXA8hxG0GgIdQX9HcB2tPH28B8rDOLhuWWD8feknQnJt9EHuLOcciM2vf/LJGRp5QikdLyoTO
HYW/UiObs8tHC75ketFb/2nOA0BltnZRpyjtP99DDyov5w1YTi6oNFQ3C52bibnOW4WZBk6KrfiC
b7SqxGF9m0XhiaCbGFsW2I1M+l7wmiJWT/xrae18N12ehW8AnNktAyZz3BWisvO9GrO3niZi0SV/
EHMiCetz7lMITq8DDwGKMLSr99e0D3Rf6+r4kfEu/w+rA4JiZ9XOaGsCBX0gbljFptE8i8PjO1PE
7No2q3PrEAaGLwkGORi9F5gbLn3rSAU4+5kD3j6+XaRSqIWzoTlny+cHX5wytf6cRcCimzVIo8Jv
h9fqgUm+xarzNBOSt9V4/Iuf2Pk0kudKLNVc2z/XvmsKvgHSEXeEqMfiGng7XVjexBVNBqa3SxEM
Oins49+vkxIG44/pTRg7A2mSfkrzY3KS+WqyEH+b3JGKg/ERo1gFCHrxFVb8Eu8Qadl4yAlV7PZr
xUZQQpi93a6zM7wcJiPzdOn7Z1cSW4ob2pAyZUj1U8WrFtpXvXsM6XTZfmxHHASZyDw+NHlMYqLH
IjZFtwn+9YJ38GTxR1CykNWWSaApNVzUMwsIqJAy6BCb9Jz0JK15C6Xyr5NNN6JSkYwC1At+yi8f
5fzc7ItCG1yLT+YGv+uyDoEBIYy95wuep8cjI1ijTySHPB4vKOMM6fpeancYWPn406fvyDNXKwyh
Teq1WWOWtrbRDpjyBvUNr94pVkHRdOYrIsyKXJwt5+xd9M2N69NTT7bxBCfl/+tg+PMZKLfwJyEy
kj0CS17lGQ8MmWjHUjhT0P3NgZ5jlpIEQRs4BViBvK/sEzXyc321fGao9hnvhPKQ3PBL7RRQXW6U
yt5JT5zeK80DXK5b7NynN+x9bLPUFKfMQud+KovTJ9/BYYeouwkvny0N1xENa2DROWFZYtZg3UdU
MKrww86EmlNa0BBF3rhwyCm64e5XFbt4wO3wFgLxFmNT62/EWOAxpENp+oLcdK1yjaHUhoxsxpU+
9gYobreisKhV+VexKdQ4yYOmdB9yZNH7XhweBtM0TBHLvUzyZwYcCEsMLuELA/HLCafUcxR5FB/a
kGSmF/dM/iDg9Su3UXW+GB3H1SwE3f5zYqnFOjQpVNqAwvfkBKlHewCtutem94Xl01WEjCA+FD+2
+89lLXprIPphzmZoT7v/qkAGCxwkRL4fLvewdChzYDcxCLO2GaDEdqDMPI+2TZJ2NX1jwdT0j00Z
MErEKFmFUYxKRE9Gx+wElNVTFnepzQOltcCZSAiOSn/AZD6z58ZWGMxl60QRO3U0Fs3gQA55O037
ilWy8QD/9bdZpPIlycibc8Vt7fVDq9j+DUQr/OdvcDOL4w4/ADoyWuUcLzzfFMRbd1cR1YSIx51P
qsivzCvh0fUK9uBUwNWyGYHBc11jqq4owc2vQhGVXr3MJReu7bCXz90uv5twpEUKz/nO5WeHkQB2
FPq13/pVxia6z86OZ5QMwh8Y+ekJsrWLX5KXZTPPvFmp5q6/TXwSrRqVZH+SvVoWjPxTCFwmF82k
DKTVZLF/UYjmG95kqzppo7xh7Onlu5OEkORGs1yWlKd3PntZ9Y95fzeFF0Srw2TxQbecR4QUTnrB
NQwu5f5U1FeLmeSUodyj8x+hUjONXGDYUGW/0ZBAxhZKqX5xWAmyf+cDMtuktGCznC4Vx/qcdtOR
Vo0miFwC8GAg5OIlF6+PcVkBg3KrJgR7Gh72lAPPVzzUqkJX8dgxeFbbsAcVYQG2qhZikHDvb/t3
2PTqGYzjJNDc2NkQp/rH3/fDiAXroRn7CMBn0w5bxungPPMUKRjdo2M37xxQ1nxNCwW38QIR0gHt
UOJ4AZ20XdFz+xW1JXbVDBwscY/CcOpB/WgHOQrmb+zXBtHAPOiXrb/YLhPeCqIZ6G8XHtsQF458
i+73/t3ySlOq1cbSqAiLp0bv1GsClkJoPO3Jwf29OTcfKijrqtdy3DoyS4+j/wFv7XO4tvtrTdSS
lLarr4DmWX5L/e6BNOfsb41TpsxsFAYhV6KrbqeNHg41o51DNTkU7b+LJJgCPZdClWPA9WLUleUK
LiHvQwE3sbW7NzTpHdawXAs+Gu3uEzuopbZG1loqOXe6VtYrwVtEWS7yvmuvZRt9LRVznsgUdKHG
D9uICJ8Hnx9W19/C2IZ5b8fapKJFltSy3HTgxSbakHT6IL68CeVmV2ISNpgjAkgKd+2IdmMkOBLl
zmzLd3CI3VovBF83h1jy26fiHUZnqZHjz/oOF8bX5g78L34evwfpjD6XlaY4NF0hXwyTx8V0hIHp
AFZPZlz7PTTwvJrW17yCZmA9Q5xqAW52XnAfUcrWu2XviQoL4SECjdo+nxynT0LWgB58O4hLoZSo
QjSB0XB4O5aQxW6pQiNQY8rQwMJZq3SxFCym/n/GiGweG0i9hFZ7LLEND2R+nTvE/5Q5DZssGdUL
XQKjlva1jRDkTxif4OnUWpfMCaVxOWgLBE57NKxudfLgpsizHGc/ONIan1UMfzy5odJ51N6HSjkp
aAs71tdfgVsbgrgFxLCfDNW4vJQgqhjSjFb62EmaPkw6IUyNqS0WWJOSMbj8AqK5XA69tj18oWjo
Y8VPoRipNVKW32hNfo5vnhEuapT7Tu0+yHOI6hQRGbAF+s7+x3YWtmfyxxJdMh2Xw4U6/bL4gDwy
R2s04v0KFHJ6HNdVYhrTb3ROsCUL9pzmXFH7At4AZJbCbyHLqgNtnP4+PaGqZjF6drd67dcSjFR4
IbzwqIQXLnCpcg6ZwvsOGdvGNe70WRZprqFDsCuKO473cO2mrw0R/qu15MvA/gK3Kix7NyX9JUba
GY3S3eEnY0Ed0EvGrlvyMPiV3fnLER6Ss8VttyLWFwa+uqxo5p+EReXEhlqNfJkWDAo1IxwuQz+B
kevgExuZ+HJAHNjVsBNpAY/kVCCIpiuhCZ0SwplLLJTa2JvYMJH/ZJfMOoXGDwO0mtlPAlnI/LCg
KLv51JHuJjJguFxL28tGveHMsuNxZOU7FuH3iDhHWkTfLwv0/c7GMcEAlNLdXqbZ5Vnt0kN27KWF
/DRWs0rQVsVX+IR5yEep/VvFgQdGsY/8FGtykKOIp5asVD91tKbZwzQLn2a2ibUyWP8XxID7g2DN
UorQr7UEUli052zcIs4fTOFSYsbl+k0jgOcq41LOr15zKsCiDQXNEVzFoAXe4LNa687bSXkwZSLi
tulRrQXFoj/X06p3dxUIwGj+wOCUFd/xubdpyPXLhNvOLKJMF3QOm39T6/d0riFBX6J4Hl+bMl+6
NEDuDMw4HiPHOtHQr27wFZ8oVWfmg/whJNn0YbhI8FR7u13znIZz51rs1wjdI3tAobTbnWM2JqCO
3+0T+KLwFan+Vanb7lQfAHX3ZVUEvjOwbog3sy+N9ar01XfPQ6uX6NVGtIw1G1nVd9QvMPO9PEmi
u3dh19yG/8ge0xtvjECdCG7yodIHQe0tlJIQxODf5J/6ffNmzcR8WfNqJCkFByEu2/bKZ/XtrkUh
PW08OJ4VP6VE5ghCttO1jHI6fMy1i1uDHlCNVskYeQiazLLX54D+G5TOzYAT5Q6XUghOD+jGZLEe
q9N0XcMVw+HOw5jwLJvDneyewqhoUlFw+TENu3BiZeQCujfXOWUJTMMZENc3gZs74byqeIhW33Y3
+6Ga7vSEH2ZeviysGcorLinHx2aQZhhArs/3BO5kaEf9ARCGcgqU/Ont7Wyxm78S3nPUWHmy+bIW
7CAY+ruoopvKhVIkq5auoRziVojRFD2Z6oqNQNSHOILDV98ThMzhsrf+2TksbV9UvTkwY2VlNqRG
Gk8jBKQGOvZ4u2IW/0zKzWQjLJUGR2pTGtaYpcOuaHkk0ZVLhnUKtjr/YuCkF5b/z9ROXq1srmMp
PFoND1ygZSAlPvTdX/ezryM6XAymp4GFPsEdKc4t2prz1w3TQLR3S91KxDNVsSsOYN6VoY4bSDKy
XGx03wV/WlgJuqpvpPuoiJF9ilQM9DYnYuJ1H/WYlViaCsTfWm1Sq4LCWqNagmzGGMLcLxzwFCzX
rx3rXgAhJD+TY6LY1aIb1WbcAinhtDT4aLgwJVe/5/usIVd5qb+/YcsduuQ92qYoDq5dqeSHcDPz
NVK0KRD4RnktyC1fzeGrz01qJ6/7WHWBfktOGTXCrOOjCMO9wKLaVdfxKVY1Onl7547qXhUeEUlt
01Y2SmCVCtr2pETB5ZvDg1wlAcT+ioWPABk/xR/O2vf409O9L6nmwDmZo4CBHI5O5IYHYjN2f5ub
SPwpZK20V/YxNzzQ+knsdXiYqOj709xlz/NpKiId1T1cNZ0EiCX/jobCAWmaU/WVXKCneU1nP/Bl
xWZiV19gD2xyP2QUjuThvhKVvinJcqYxDXRqgR/r07bK2tnbQo14wfKiLWXh2MaiMdCWJl6nVaLU
0oyWlpUAsTII8zx46hQbVE9onZGc9n/ORLW/hE0a0PGRIbd6TSfL7dON4/GLXM+3TbEulGUTb1L3
GHhZwR0m+4rr0bbVjPAW8udi3qS9RuntqAAS0RunRO6Fh4ogiXijtTu1i5A5a7SmF2GGzXnMdZWl
wn0DHldqpZVP+9QbwjTAmQbAQ1/3iy0tPKV+MFK5NFfwKprxffSHc/+Tci2yWJoLW5B7K6FpFO1p
TfZUgWrY4zOMax9eWs7St0JYJ/54laDTTYG/00MbkCaDrbyhpxEfHqSaTiZmRihgMJ6YCzvfkHbc
2t1d7aYH+jcjCcgajUL/kXvTEHnSPPmFaKk4WiEJEaP3Cz4JZkbI601oEWbvlPhy8/rA/25sOj38
0nNjClNNbNjYLLiAG+arKr8EgWNTucO4Uez6Kou/hS2P65ZyW6LlFK2qbNYd+2iLZhmZ8k+v1hxj
sgiBhh+CY3G+6TvNaZ+igt6e8I9MDPgTy/iMApEtBPNZ5wfjucxND1YI9qfzftRMFulRVen1KDaf
rZRATrZEmpTBms9D8CFPT1hwOL372c4mY5vCR3/Rkjp8fQkN/mtUKN4uqOkY48ToRDYZURqiNnHA
Rg5Eoxbaj73uEi1oNpuuI/SiWUW4VWaleGX4pfjK3CYLaapYCgAl5Mu70djNfOxhatRZd2ArUoVX
EHp3IiVdNZ98eofZw3gN/M8vFC0cmypygMNa2cnOephdMMGjk3AERJv5kdEltTdF0j/cpV/POw9s
zJdTjqoJjOkKA5sI8KYiK0fEVxOIWArkLGKhFUlBLGF6Ruqqi2IR3QcrEqel+SCi90jMfwQ6XcQP
Cam4xd29rk98PnMXwqWosNTJ8ZWMvGLwfTUGfu59q6sk/zo5QA4LQivtBHiULN+Uor0lawmwwglR
If+j0FRc5JdmKUDpkbSEf8ztmbspYqE3ARlQJ718LBgXxjAqUTG9pbv0cpmA5N6aFTam1uufdhZq
fFdp9gvMmdejZeVpiys36svBFbxa1TfJEfsTgtXyeH387rMzRXY9AnlAGB07YWzm8W4CH87W44VA
ff1j6CtffsTTXIUX6VZ1M3ehCAXoVcgre/9pMs73/jfJyMLX0yO8X8BLAXn4n0CNUOEixvg4FWtE
ksZxDJE5dSDCodlptZJUKuGn5ysUptmnn5xI2Ntq8ujSzo9vS/KgTIXX/GElWWdYftCpGe3Gr9lk
ixcita0Lhzm808tsTr2DtepH09CoagpMuxM8zOWUt2a5ZS/GKNETp39GQJCBHlr5dTR3y/+qmWid
dy5ekdPrxxDaoWXdvNojyj5xwZsHhalNArpJYeIJGE639lAvx+PbvjWRrhDi/gzSGV8iv5LQ0CQL
/cghk2vIZVN4iLjYprVEhCBsWLnDpNbxpdEpODr/Hx+PKW8wvdSWH/JAddIMVt3tnH64Mc3nKpnv
wYFGsy8xyAh9NtYp1vwM9CGUASs1EmPV2/v74blqnLar68LtNQ1lwNvfu2Vmg97GFgQ90sv1+DY6
nL9h/4jKTnoyVJ8Ym0AqGNyhDElNPZH27dsbbWfV4kyrAJ5wh9EPkGVTpL1yzP+wFfx2HEq0WEg4
8orGypGd1epAJtY/Iq8vv43R8m6TWmsmRvaEq+oW14z1SmWjMfgzl+Ztz8b5KjiL8vpJ6pCRhxis
TOI2u+Pvkgd05/eyXVo73VEwrUVeIpT8rBwz/gbECfXfDAC1p3GDU3eOO60k3LaHKQeFYCogtzTm
KtJVxiZ9NrzsR3i0uuS1rMupEyKLJcnLid3HpHJ1RgL4k7q/oJ392EjwPGqvpibHinKUl7eeZoS4
n6XW6yWEHFt6KJGb0G7tW50vGJds0z3Aw6BWBCGMFzCevKJY+uG+EqqsRz4McgZDt4UrL973LTtP
zq+o/uUz9zctxDG5irreGoPGoYboifYjf8GeFAZjY7tDgdnTDw7R6gEgRMVqqNjogGlqeVltqIfn
n+40JjHNBXwj55jnWLkpXhjyChhGFMFPU4HzZ0qa0z5gUg15JNA+Ns3Co1CpiRpOfL70CcAwYKLS
KGgnuVgTkCO0O9TbN0ijUOrZTQRrkoHTpsFI/4qEOhwY5t5DQYuZEdCbvZw4vnmkAh4JydhtDHUN
5ZCUQtXMRzLYo41bX6udwmoVMwpuJBhgUXTfN+ws0dAQ2K0l76W2/QrwWg1p0GGtIVVPTWQlgqhz
9BFfPEbzhPDqYl8loCuuOILjpAiypVJL3jcLvz59dahCbZuaUWVN1h/sBGdNu7gxitMB7CrJyN3J
BzGnkEHES9sDKlndiy+xMfop0GdBqnmrpSgA9HWOGlAO3EiUl1F3qR18A0/OUhUTD8bleWD3WGvo
4oqftVP26EqI28KXBwv52o/5ch7nLxoqGyMtyfPF2SJp3VJ427nl/JSbsFoDhe9amt5PETt36H7T
yY9dFpelK2rPfhi8czi35OWHCrba2OWK0mUDiIo/v6PaQcni40l70FTFAr0ewJWBYgkQzYWVNxxd
EaoJ663E6cml7WLwuUWseAWkJwJPXqeJCxcrlAEsKhrwD1GPkqfImyGxIKJE1ubJ4k5oJzzVBLXe
Rv5Nc60C1wL1BD4W4MvgWsYZT6UvX3I9Xupac2nK6JIn5a3utLZY06pnI2pVVDwmlsfcJLeoH8u6
Rd3N7NbmJTh6UVaSzi4wa6MiiV6Ij0AmDkCk50Mfl68sefP9uNBqD5KHYv4fSXNV2wQgGYtyXOtf
hDCNb5NUqe9oxTfhzfeuBF9jBnV8b6w5WFfAkXKIMmbSEeOSNcg8DoQTBP6QipCuCf5WN9xVWUhu
a0IFzOnnMxmQhDtg0DU+3TLTdiuYr7YZXlY6ASkAeALCGQIDdF53mndTZblHSnN6vJGoI9OQAf9e
5JoU9+pZMRL8xneW5xoPm5dTTXYil2QnrmwfwemtULnosmVd11eGNkfaOKySI2AjYKKgO0z0JX6G
4/WBhbVh5qgu9kxFbWRR7IRG+9u7gIiIAolFvYGslRUNNUQ9wfP0EQV3/ZuzremMOuCYJ5cjOnIg
QwLuSRRr1t1ry8DL/hmFTRuZIX2VRj0DIpSLxqGLSTR91Atfg9pkbibl26bO4KnZyVdunbKXTCYJ
ckvvWXeqYrAFyH6v7eqRu/Oir4ivOkmVZBYE0zanYCA79PKxN4Wk+0UturQy6tUgwtViLq/l438d
JfAlc2zliK/s3Nc/KSfSx0e5bN1B8FmQvunQb27jHw+VGc0y1FMiY/kkI0KoC0hHT/6CZ02iC5m/
Iylxme208i0vThkkbnMd4govLqKNEB30CtLhpv1+UeR19gX1Mbc2Mp93Jest3bH23pzYlIHulU6C
SDZekEnOmV0wtjAa4HRWBpIAjZSQx0Kn+ugfQuRY5c7LEPpIJjXSJD8vF47qA8/A1Qvx8x2gGalT
kynECWKElv9g270JVXlsD2g7f5qsEJjxxvXOfcUIOz0LPqfrFIVtphc8BilLMw46gwcTVU5SxMoX
g1QclTIAR3R4WHfIxIJRqMmgitjahwpX5SV1xzJk7omGYkaxCKUBJ2uIQVAwqihRDKtmFmmpuhOG
tnegQoxqStmYq8I6rFbpLzPNaT7eHUq8QWd/98xFe7j54HlyhIlRfSpAxBxCqHzdE9Oa3tlBuEM6
3/1nQutVi5iZYEK2gTkNDWywS5zPqDLEGLbLOwEMnDsthBtnousyy/KQLAvPevWtGq7d2YsnLZ0z
Gp166g+Ph6mTFqVgVVLn4F8eycgLyFHkABMTA2sxquXJW+oH5zGJRIbwOEVm8eUUaEPNZrZObDT5
sUjFHDhfNQTDSdKCgqLDm/+xtSI/RM0UWniijhZ3gZByIg96h5c75CYsiNR3z4zKtyZfeJVu27/p
J7phrI6wLm1eF1byhQHW4vgVH8rXicHYpsNiPqeyi7aPvh/L4oG/WoUyw/xHI6CdXp/gsWrahbMB
3PKrCSFd0pd4mKiAqpz3xqnAwK8mD7EVHr4RxQ8qVA+58Yi8Dg7S6g2rpJOcnb+JWKgUntiG8udb
L52u3jdfYC0UCEArNV/tJMATQPQg68O/e5HmbUWGLtCHO2f9+diRfJ2Zss6Ec1nH0HMM+MbcINYa
t0dyq9XYvrIXLOEMOZdPJN8SdvRFpgHRDi+8CC+5LtqIAgWqIT+W7XzeYh4OoXsmOvj0y22zygXa
nPB4wkdUQjX0ZyEL+GKdZ2xie/+7KGhUIyw39WK2LVFBAd7QTdKOaRgTgJcGTSkAxRcodc+Bz/TA
fjcg6+eBwZb9oAzrtF4mqJ5YISzKcGDNSNCEjzP8h7xTpjECcMiCLd+xJMQaLRBo0hDXBJ+av49L
nUCDckUQWoISkEIZgUtbob+dPO2KzW1K3uKWSMe41wnXa7SpAD2LNlCkk4tSNrQGvpxCfcMnl+Z/
nI+rx6c3SEUqLUtsXOplr4ZoZVo1+py6L5uDHQjdQRtbv+HSH9JSlA+3MLH6e6ign/CUiRfb+xgI
+2YzHeeNPUrnyi6ARoH2L1UFrysvtg1oLgGf+Z1rxP91uFMGLMe02HYqohSsJ/l09hj75EfASnYO
VPTJc0x/tu4GeDoNZHRiDq/HPP5cZ8aT6Fy8xZUkJRk7Sl+2yTYwla8mI7qmDQGiU8y0TL7pD8hU
nrYipLJkooC1cyZdlI04izFrOwvFl9uVEBNP136nySvP+3YH08ZUrwTKznnZ1+/9FhNgiSHK06Ty
N+NFxQ+r4Twl/idpq1ze4JW5p4AFZVPjNBxC9s9pKVpw0Eu5zLGXWhECW9fvZ9b9V+Y+fjYG0d+b
xRHfQ0EzZGRMBZWhhsYqKnRNqI+G43KgB3T3B+sUSmNOCeNMaehj6I7Omgv5LtX5q77YkykLGjP7
ubpkPhZiakY1bK3/9cpx5SKZBdRn7UnDePZTgt3Zi1PAsHblcRbApCdlV6drbv2f8y74r/pF2Atq
VIXdKU9rRiqmFjT+IwjoIb9YyCQOv4J/0m1Xg6UYohxnwosA2aS6KN+TArRW4QnqkPoLtm7j4Vq+
dtb3UsgZFstynVEnQjDL6FAcTp4OrFQmPkB7VakIXnDd7qTyp6VFBUw66prPxNpAw66PNxWa+BO3
V5Hd378Od2G+nfEC8/JXQxK6h9+uzHrGT4gtqWxuAoQHvcsLkdG4DZdibAOmPJTPvrr0MuwEkUX5
VDDRZopwSHyCjCA1EoC/CVyWlhdK7cOoOchUD8wm4tds768Nswj9x14425F9aIXWJDEOniXA1TR0
HpQDR4KGa8mugtX4RJLRqTgNuiNZkdLncDzi7FRCMFa7xh3U36e6CQWdPTW5ZxO3x9uGogvmO1uy
mssgNnFuor+xetwMNjq0pF7YHK9H2hUYnjK+fisFksho/fyGc7I5dheg8yMlhN3PGYuJSmGUQjZu
bvG2IzoS9V4qwgLFZdsgf+2NQF2bDR7xmRh81rEmBwb/GJfk0+C3T56rNRSJ3e/+1iDU2aV+4Anz
4GL16Uy0VOMnYFJO+mIQEFQgusJeZCV749Tgr6vepbFKBq8iIu8sa9H6vDlDR/RQ5in1nj0lOSeg
XykvkzHE4PoToF94qJQu2mU9h/yU1oem0quO7lZ6bEEJBtz2+9z/OLAsXje6M9Qn6emFJx7i9tS3
2UUDVyvKdyNkdKoKFqOUO9YhKOWu9TeFMdokUXkhIB6I9sVoQXfByAUe5B+26hLU1uWtvSbt7ewK
W/2bzwxmN6CHehI9sezJDMPLhrxml+ZiDugfIDEiUytXAWyT0Zw9JK6WGZMUUJMDe1Rjvs4KA/WL
SLm86HPig0jBjLSPHI3w+60kDi3+wcmbFG64HoqUtyGKjjYGCAfQ7Fh35dRjN1uGmn2FBB8gcGVJ
GCRU+fy24TznwwJ0urMnbKhWxZOMxf0XC/J/j4KP36sNhfReLJ8g2Jfc+6ve0c2iPjWqhXvrgsiu
3NTDBEyRbt7N2eBYo3cMfELhrBTlP9rimvcsKMc196hy02Wkv+JmP94PS6ohBjJ+icxkqtKFgvTb
fO0GBY1f2igZ5UCWL8NhD6918oYS/RDoFA89joAUQdm+kAqGF8qDJQ6QqGjRFcWuWXWfNx9l6fSR
6g1lB1ZbBAyen7z30HAjOx1hU1W6O+tpTXfDqISgywBjHJgDwBadH0oN8Oze6NpKjhlwuLO9yxHT
ZIq/DxUogkw638S/P5vrCNzvuOufyFCrvoMCrDgv3zFY+VMvqfYltACL1ij+mbA4MsZAl5pTn6nh
0Yuq4T5s0ybI+zWHNxdD6wuFCbjbI2RXuE5sK3G6pT5p2hw9wjBUXpFUDKz+stRKisjI3iME/tMc
NDBdDPa2lZIwZo4OWPbZBEbbdCytHzcnQholqFWgh9DbyV9zZfomdxG21nNGTIPIi7+v83LzcqZx
DQThXDrhYTzKT5oPvgghW1Xf6B1B0UnGwRInbvfQxgEDETh/Dd7z8e7pl5jvTlsb/c+rfxoZqv/q
0C55jv/tR2AdxUoBzsfYe4q2RZfk5fqSyjdf+lMDyr70/oXibNmRbfmTFJJlitOgTa9ugOGx5JLZ
zEb9sEH2+J+cGoCtiBrpi98onpKU7jKxG+2ClGnmqoNfn1X0DRACLI95aQj0/sIZKpsg9k5f0GLI
uZlCehGrE0h9GcLTdByfVql52asnPQtfikU2YO754TYyujUPXi04KiHfj2PzyGYePcp3EVQjsFFl
vtHLxuJ5wRkTRZ3JeVl+cimGNkXFofEWTwsklB26RIMZBJ2aJDTGdXTQ3lP6l5o0BkM9uQB2qodv
RNYeelTbNnoL0oaRghtzFetnLB+bhrCzqaKMdEZe+H0AnWrEkJhAZXJq6cNzMMgvVzczle4L/YuB
SVmP/cb6Bl1a6e632zxJR68BgrDckFnXrS/XjGAGSnREJTGc0/M0OF03M3xllSGr5wo+MUXzWZYV
7FfCt0FgR6ldcEYPhh5+cOiGWcZ7v1oudnBAg3YGTled/Gld76AV2VGJPrLrlRy2+A/t6Hm72fAg
LP6uwLF/exB0YsmKAAkIROmM7shz+hzsX0lXT6I7SHKKLG+QPokc1H8nvlK96HzlUXAfSA1grDNW
2vn4KASuIzt+mFlmOkR/Zv2ruSYsqRRM0yKhylXbDKZsgY0syNqwssDqc0d8WyvNrX3jJu571pGt
KKUh2weIzKQF2LTBRgz+K29a2HuE7JMs8RWeWzbVImtBAO428SpIkv53uXODJQM9fOyHxw5qoRAy
snrnfzcYyBo/WfHjxt9AvJz8EEiy8miuVBwtlUzKrduBCuiD7bOkL4OKf2a4dsXXshgDAwVOL3Xu
z3uue1rW7jg9OxHJZVksA9GtboG0gfTRm/CvyINsc/Oc+kmjqQDp4GVO8fHgMiHrAJ8mLtqLHOo+
sD17SWbXSJm8ryhR5ycxvP/qveTb+EO/zbbJ6BwroiSAyFuMdNxSXJRNo4+eKkKd4HZTWFeZbkpy
TtOX1LQpm3rtM6JGK0jwXnN7QBFG8jLBkAKGoc9UUwlUILrTBfYeeWtks0jwcHH0OsUiGIviGyOD
n5maawgllSgf/JtGk11LztZuY6L9sn/jc7/NFGLT+XC/yd3ugvTNmlRWoyacHl/15/TLefvqPf7V
VOBHDPxNxGq4/Vdve6yUnDEF4BcqvVHdDf88Bp9K4TzNZmmMvd1dpxBR2G/sK88aQA7gHURrHB/6
BxK/XEDVD+FVFC7oMb9sPw1lgRZJiCj16cWxgg6hd1kgLGs5gVCq3k835OqDWLgwdYQ1sUp12Rol
+tGfiolpqsHmxNlj9lr95DDLlGVqOJ5YnPGHoiJZ4JufOlc3H69Cjqmsnp9qDNybY3K4Jhl2L64i
X8c1amjcxoby4oGQwUg8Ygo9eWl2wxDxou/UaaQhxnEEAODIanF24Sne2HIoTCMOxQ0RoV/v3ObM
HvcUjAsdOUcvavPER8oMeHNIB36HPmKVqKd07PpPGjxA5r0P3d0Gy5RZMvFUw0O5x+zcLYMKRUw4
dRY+GOv6OevfUWUO4RVYMw3t3ukcuDWUxdOZuIj3gECmcyQfR3dsWoC2iMSPDk1ObeeVGkNYJ+o7
JkmhTHp7N/JlA3IkQHNaZIYgdvWYg5eF6twdxx90NQ0l+bGpUtvUF3jYk1tTVFgs4DtzBlIsfPLZ
g2Eoh+Qbyy+hGMuqaU9L8JZXFszxn1GSqoePlyMmtNST3ZgkKoxZKHWyYEi9Qf89OXbz1IlIUNnR
OxdCzP4UawHnuStezstNLTft0aiQRwTiz3qEKB4jBlEOmzrZOKfAjonus5FiT19+1mep+EKkNGLf
70SuhW1GFPmgdhLVXXRtDG+kW4h61WT1PhafNzOdR0TPXrvS8vnKeyEjqMnkh9ape2WPS0QlvVa8
4TCy8FkNqGD7X8QlsYuBupU3UkQ41GcS1ME9PxxVYqhOn7+giIJRpqq8BPbIONj9kiBlQeFMSSvO
ldWjPAxbjMhVcBwALdM1doizrp0+vT40aaEzuh7h3Uz4Gcv/I1j2Umq12MQGIebnRWs/dvtBuBMJ
1mDlX5ByYM1P8gUxp8jCWZWRzy+4BxxqlQHaJfL4m37TX1wylHbiVf0U1YhoLVQhIK+yrXn1A7N9
Qmv6W9MdDqPxVRwebUhq50v8+wsfGip+LaskwtLF/L+2Hz0AnrAY92ycN0t/kqyoTEKeGYDTe6Pb
FOsUovXB9hDPKd3JnoxL23cfXeXzUFTbMGqSjRJOiRcKWLWmuT0hYCfhMotfaHgtd3XoIDhobCzq
RNa5kboWJgf9Nmmua7nxHONtFVP87JHHjYHR9G14amJybQK8BX7GQeWAeJXGn+d6IPg4e7v0T0j0
vAiLUD35/IjrK1ny1KmyAqO3kSsoMS1gaWPR3Pb1cE66XRl/jO/Evwr8GP1f0WarwzvH92MrQj3f
UM6TMjKoeDK00/V9uRoVqVtkVVU90PzXuKa5dR53nbatUaV4jOP5YfGDWyRS6KVTrbv3WW51QO0U
a72hYS79dK15dINlRrr0VbThMAEEkPtRLfH/XZdA3DZWdc1tEc/26iis/5YFyXr07BQnkOKYgm5h
YA2Lo2N5ql9t0MB1IoMjKzTLkwUemoDqL1jUKe5WCczWDgY/KAUwt2ev9reqjhd3xMWRgeS7VIiP
mMG1WTyBh2yS0s5HM71lGhgSF0lMP3lt+b2AtZ0rT7F74LiInfuH/MlfW2i4gI5OkoR5vwb06rWF
9OX253ElilNbqdv8bmdBP0edKRciJh7TcPSU+05T7YkHdCd5IK2dMJ+fXu2KZlSSaYG3Irdvfrfq
M9p04Ymkm6p6MsPIOWSqC/4VPdZknCB+ylt0sn/VMTj1b/4vxorubGUHPxvQpHcuSd+7SzgtDVBM
uSdQxeIYbekT7+LxHatuUVzG/stY2pFeSVB/RNGvGAptK4ixZKhaYZbq1hfFiLKA7V0Vweb1Zf0i
5Qzg9KaEBvcJvgVg+3qLhMbwYk2fo7KY5E5RJQ06RA1nlT44FOCemQnNSjnqe/BORuG5AwuzmTyF
9bH9+a8y12I3S1/bSZzhNDddTNC5/jI1iRmlj2Uh60R2kpKLhM2my5XKpK4VKm5Aiu642p9hnY3s
Y5rbXXC2eU0hsNiuxT8xTsaSUNQr51mAkoxLHlWdWk7jBH25qztwDaLbcvkDbk5JtRHozI5PzPeE
cmVVkEhaUj7qEg6YWX3hxX0GF3d0bi3ITHDeqQ8OIgI0ZIxvXw6vfNYA7ofosvj1zSbRFggdrIVX
EGv2BpRYoAj+b4txcvdezIgq5pu1kEpSrWIBilkREBNUv7knfXfaG57+2t6jjh+l0XOa2xwOS88T
6e9CDka1WBFvpPBE+XkrnbxG/yoNesI6tKTwQoOe1oFMxNlpMBivL8EyWICm1NeN7xpq02Je00w2
7AzLKCZ+a5a7OUuc6PoHigcWEnkasENvyoRbHAgaqAdDd1lDLOfctbn2PDfQqU19vL86gcYCz1jR
FeN4YfAg0KgAEHVpN5/W5io7H+2ICx6csMHaHg8VBKc+zrrN6M+cuP86fEvrNuUckl1kMJ2eGR6g
+jDz6aM9hlH2yZzCLpyEakie/pdY7yQP+ikqyxPETdzU6ytP6cadeKKLtlsuWTRhoBxGTgyZqq2f
YeFibL/cqJ70MSPErKXRj9lBMHCVYjMyzc1U8n7NO7t42rNrrb/oz6m9nVEe1g9auZPQRop4OE8L
wWMncnwTp53Z2GOdFfAK74veOQmRDWMYeVINxv0ALi4NGwWRTKfiya3iiEfhodimEznUEiEvGXNH
YovfuQwwvpia27dcQPmgclTgQ05XVvSXcBgMFq8sP4D7Ja1a/1GJx5IXLujyM09JMqFTuMgRcPaL
zYKefS3xKirBHANmX+A3jrydwL4+52i5Tc5ACMnDYpmLIOVm1HPCyBFwm93u848eFEit4AL7OelU
+KNYMzIhAhQbeC4xeABkpe7CmIbSGQA8/NbcM2nHIg2xV5odJULV2kfoql3blZLUbcNTfsI8c3rS
vH69uFGxFGHWsgIFJvBybcsjhcxFH0zA/rRGKWnHfVz6L4bPrnO7tlCOGZYc/GGdf16HeugoEbII
ivitN5kJp4/DIGhjeekI+bl70ImhMw4+31YfNcnRdIB1kOLFaLc77Bx6uJWs47LAHMzgh945sgCd
scjxtJvN3cQ9KEGQHIbJ7dtd3e3X5zDGMT5zmIPut+akpkPEU/pZfQNyu5O6sN71ysZGDZIp+rgR
tZ7jFzSAVpJ6oJ7kAq89lNr9dxB6urHYfpEupgiDhwzgd8U9yxFM4mnqg73EH6yKcj5+gI8Bu2hg
xEV35aEzqVC7nwgqQFmNsjFA7GnU0Jri74W3HcW19vXUaRAyBr8vSR/0ooNhjwaXoJGtxZ8XWPu9
MUTgVjBO/PZvmi8+qG3i9xIPeU6ete9PSy6WoWGDwItIbhRWkdiM8M1/ThnLO8EkFA5iEuwWPrwl
qEUsUCY7rDI9uCDhEnEBOq0jyLhtYBdQ1rWTiE92Ha/iECJ0Bnzb5sw2yHewYf7JzIU1nF8Mr+zi
Emd2RJ27V9E6g8eALWRl9272NpZbbrdtjIMH2wp5z355mms4rt3iOF4cCvmcJJGK8Fkb7IKubMWb
DuJTNH1usbigsQp2QdzzakhqgQyG0J5vdf9TwiHpNMN4lKG2oRTLDRElx51rIgTzUm2Kpgb/RRnY
JGh0exUdUnIhq0KTiYNidP8TjanYoAwy+LdfzYQ48EbC/iKXbTDNuAde02dfvMhZJ58BNu5T/ugo
/v8acWKbD31NoNqT7vzWBAyZ8d2WMluiGpC57BienqifBPrNk4w8rs2UKdx/fMWspl3TRJpeAsMg
iMXGBfA7+9yx2GscPUOsWfdfQwNoZ8CaUY5RIPzluK21ZTeJ9j4J4xhMn4iheKB6X149v/0oOewr
cO/hXkNFkHrX9IWA4NY4l6hmCtPZK1x388NB/3sFXIVxksk960NGx9lMaqCa5xY1Pj9Bl05ck42S
p2pPTCmQWS/SXifG/A2pZLSM75hF9JmxzkanMMoYDdWw9V4FeU2iDlFppbxzIgMRFbBXVsFXOyMW
+ZLN0t+4YWAaM+tAd1zHAfvFRICvIIJZWpVOQhYKqLV8n5Eh9pynUeYXRTfWpcaFww40/HPKSZc5
fR2YMEsPDwt5DmviXTLM+E/VhNPqhzJAe9RtDh+ehvBI7AxucgerXpno//NQNg2i14OI/Bsgqhoa
S1uhYl0TFjkqMZeGcmloCmUMboOCQPC3vCFw8lG2ANIbMDpzGz0ZRsSJzA1WB/y58vLb9ykhBpDr
pbodKvoUqKr3x5XmEdR/wUKpxUaWKAo3HvEOgvg6IS57z3/GPKBhjcYljLWpYE9Z1PLi4D1Fwsrk
QfiBB+Xsj5W9AYhKAUMMhUktwR/scc/YJ2Rdykl2cg7VsBZm/mdR50Lv2IlV9IciPB7jQJr6jbe4
8fkas0dVnzSA4+5NADl3G+woR1h3RGq6Unvt4FH0pVwseKhPjWxcmj9nG8O/QdBecTUHb1Mb5D9a
yBCPyIfaL6htV6yE9Gh83O1NrgDBsPtz5yblNgsntmykMFNv1Azx9R8mxgN8IO21NnVgA6ojUYMD
UxfjygivbDRY02dC5ioFfCAbbss27tbXnth3gQOhTCj9TB7OGsvffr+OULFXAAY1lcL+t2Zh31HR
ik5BrIbQ3tfxjrVk0fdfGFFie4JoQU8Q3ZOdK5j+aChiG0t/MGtj8E7aKOq7/sJcZi+Wmd10Jjk/
qJoIeVrLCoHNbJp49t4kcNj0AvP6IbCZ/rHbAwpUoJ0VnjWlQSQteVNS3VsnSZDOfoczEUo8oEde
7HKEwk5X9+05t758NsrLup/Fjp/wM9+FKttjtwvt4fFNGHUyQ8eqmuLCXK/InvnhwEsW0G/8Gbp2
G1dmEqd2jvxD4YwY/675IEd9Nla9Yd2K0LMhQJkHgq8ilmGuMertt2QstXSogKoJdyKPXmjm8w1N
2c2B7f55FE67STHJDTumTESQqhvzdNUZvqFUpbq6T8lT7ksE6MA2Ibs5csdOCX9XHr/bNFYGaiNH
M2nRDsXdMwawrG8qsQ6dYUc3+vNgpa+DCDhaYbXV69VQkf0vUELPYO/0gqsRi7CRiWCyxcSJ2wwD
5gSeyqnoqGPq/2BgSs10ZiREvwe7/YOYyLklqStb/pfiU4YQ5h7VDN9WiyUreVXGCy+OP7YvRU0d
0gxaC3cQK+HDeB0EHLSZJ3sIu4ZRXfHRTBaHomP7vwXHHADyh0GuJvOar8sixYlKbpq0ZODpt8r7
gqmyIBeaN4juP3H1QwLmXjQwWRandlaH9L3Oj29l0lwU28RlpMX7U4g+rqVQOqBBoyorpoynrrDo
lw6cF5/6vG5t63Xeyhk9gQ6Dq8Q+rhEbN1np0i9wlNW3nsUZ2tV4NHAVp5FBCMoZAiynrI1/XWQ5
lTl5zxY3S50cOUciPgDeyFbSj6tUUSjkaSyVkWDlhddB+6s+ZKxZWywtT0WfshTCB2UeVTqbjE3J
0bIdDPo7aHjnUNULS+J8nFItXl9XAQW63dcOMzDbbpvGfko/DPgoH2UKrFzHVGvpde60p3x4ZjeN
kYXqg/0izGYgS76VOLK75yKWtcgMQePaz82Q/5ZpYcsQa/QjOBRAvgOwc3PGnXb+a25uPVFy0Hum
GFgUlVlbjZJLXFm10dI6Lf0UDxiFWZS+NwX7PzijyK4iT4XFd82ekO6ybj1YmgBVBmzOlLEngvds
h58XIT5bqNGck+cD7UwQbYtbfaoPWfMHVQWAnzHHTfuZ11Uz5I0pLW1parTvb+J7t8LoFu/epsDr
V7e/dBEaIJDfJg+VO/mxizE2VLASRfqfJWc0w+ZDa94FfvEknpWXVGd/Sfl1R09B881etfYxhWSI
LX3Pb5GcPAzYS2fVC9ZAnEAHk13xVHAjyQcZRBVOjPmzhvjIuPOd0trB3broo82FdOMdpQmbxTvH
oLRyeXJdwsd4S1Ac8Xr72ssVTY4zlTp4Bzb4Ep2peg7r0DWp8wd9dqStQopEX1Won8zL/qJqxQSm
Z4w+pUz/VzWXFtaOBtAN+dMN/0KH6jGyhD5r6mPu/p2uCwGyxPoIBeHfrw2z+Gc+0OuGdMggNali
o/0HCI2WP0RfdurROiifwmUbbPe3mvjIZHSdhHXNYogQNb9EJfRBktvoHmS4fK2qHtgmECLgudoe
1k/Df4Y1IKmOcmyl6Sv0alP6YrM/sY81mSrwP5KIMFMUmejX9d2Oci9dp7MVcqr6y26o8RsJ27+n
C7Wd1eyBEIcnAF4d91WgDqSxAVbJBEMZ8Guv8uU3QGknk/ZychVSSnLPhKs9hyP4xNa6RHogvE/g
mTUiqNcohJgtvFQ/a/tjqy4dR69rOCzIsSqMAB9qNdNSeeUrxcDeGPsIjjtX0KoeTlQyyZ8WEb+q
tY88QS4xdXxmgJjvdF9v4tW1/M3D9i35w6uJn6c9fmfyVmSOzKHW1EXfnvZaHWZn3sSdiu6gnzX5
UxGMQdqHgZnmNi1do5GkCN9tuFCG2K/onNTkOAulAOVpDX5GD3wFIzCf3fFEmXY23dx8PlgDW7xJ
CNCqiOsO9xSp7nJMzvN+d/ibwZyHSyEQDpnSKjak3jobMu6PI9REQ7jXHpmYZvQFBqU1DbHEsKPr
suKgLF7QUhSRuJX4ghDhU78EKG77VFq0mV6wRQjgtVfsfqmGhRX9QYaHj99TPjcJsfGTOtnMqsjV
jIPnDnivE6YCuKZQzvtM5Kae7/SyxJffhdKblF0N+oztwB4SRxFJGEy/k5MkDj65I4r+I8ar/9v0
nxMbU5RkYNLretFJfNp09dvWI/VAxOIS9yyEcP6PmzonJKOzBZFME8e8ksAFsnZ/F3goIMMWq1kL
uMthDvrw2C8K3VWCPHeEy+wje6nSIsTsSoFtFwY05gCSTm51nmPefv7jNOiOyxze2jsnzCIffTFY
fvoTO6GgOe9vcjTRSoW7r0wVyZSHgaZE6tBNzs2KJAp394m+YJNB1a+R/hz7SYG+/lRDpabJzm7O
/WiBn45IHM4YGhGZfq98zi51xxOF7m+AJu8TiaL6/pNhlCJw+MW1KRpXwzyIh04Y4wCXG/Eugq7l
YmWwRxUtzjvonC7tzUyT0oyklGYSu1kGxe+Zpkvf9YQPGDFIBr6qR2VhripKrYxa9WoSwNeUxHNu
VPIroZ+XZMVSxQ3Kje2Q8j9kzp/iUNkuTB0LPAfbzTnHMnmTzCpKvgM8Rate94iDZ0y0+eszTien
pkguVDSoJq4bQ874CoKKbtXSi/OibVl9W5TsOx57dBn/hxRFo06V5j5HOxxteAtTi4nOqsrcomzH
2gwn5CVyXQthGHIrv9nt9mhHZ/QQ+zBFyfqsiycs1rc2qDN0YhzY4eLXP18bRp8GEBnD/vl3yRG1
66Adhji97P78aGQ5DGo+cV/R4xFhnZ7FmkpDpjnmZdqoMyj8DqsJ+OFAOtB32xe6Qn0b5E9VcdIv
8OmF49fXZGL7ZNRfgxnPVyaBLbx02RdDOZE1N6/07ilAQyO28UsjlPec0nb7iPm0janIKYcdNdmp
pcxxl3NOImUHmrFqdXYlMNdwEHDjRi8UZhjRKa4s1vku3BBMtnr3xNnADG6le2eWFdwqz8mfA9tZ
DQh7Vt8p6BNdXt6L4Sw0/+vXt0u6R8bMDRodAjiL100gqr5n+VGIA64lbnzhGAfSm/PQSH2DNyxq
ZHB9ZrCGNLwJy1HJ9XuXtAyOa6P6vrnU2Q8pVuE+s/lVjejk9gOJZvImHNs0s3D1r6aydTBxg0xz
5KrJFynlDHo3SwizcGElT1MnFl4M0xTAvYqXyp5qGioTxkTfshWh8CDeOlWDDXfJYoavik+Ayl7z
5+HALPKW32bzfSQKXENZl+HwT3ojuRAP9/nfKJruKKikQXWa5hWVMQ0iraJCEeJc1T/UJMlKgrsn
sn6g/lV+Zo4DpHcBp9JWJYAy8V1NQ+g8a9uDOiu8ErmcqtCm+2p4PN0l+0fu43ol8ingCLI3FGf+
EF+iiKR0q1FoGL60ZcLsAnpL4ZfDTSXCy6aDStGCWxS37wo9ytlfE+VV1W90eWy8MVCxoL4c6neu
A8v/Wi9HK3QIq93syupl7z5fSONM3OhaR+DcDyg5uIK0igqRChqhq6RXeePMJXIAusZbCGv3JMBi
nLnl5v/TiJ7QZomUk/mbzKHOQAa7IeXPQ3v35W9fTU8UDKu9avZyRt75P07TGv6ZZn64FzL9syGA
PlvaKhzofFt2ebLyJuG2PBU9oHPnVzvtEHf+RyYIRhZoMCYsnstdQ5fYE56bik0cEF8BHOgPxZxn
gAz9S7DnNNjFHX2bUip55V7ARc7LKbBlWWBwiwlZTec7M9Uhe6NlZQ3PsQBZAf3BAmJ4c0s6RgQF
iN1B7A6E4AzIHjjSqROwBzsNAG/w6wHjs5sFsLPxSyIR10XCseowiJ93n0/AGhziPzYBektk3CF/
Xrw/K7vbdcWpk3IGQ6ltbqaUoBHqwtdpk/S1YqjemulaLqZFrclBewWPboqMQtCjiURHGd0QrLGA
1O2JSAKAvT4fJf42c4rmd4N+HdKnIR+MAoof4XOlopoQMK7nxaOYYEOnqv0W5KstHYoCz8HM5FV6
ctSOS10+2X7SVR4Sr9ORzaN4XSVv/x5cY/G8cfiZPCtXXo3ovNA8EY287W8SZwpRxwW8gvCexJYg
/0ASCmHNmIejSF8Ju49J31HK7WbG37TIHuMflnSJR2/z/d9MLFinuaHfLpEy0IIIr7Z545bzjsRi
PChMhuG+77/vri3Ea9aLKYS42t81jIr7xIyKuO9kjV9/OwKUys+3R2lye8Mz8raLicFX9VZVAr4F
l4mAI1UwXNGJ/KrfExKnb5DavMKUHuEKM4P9yscN+mA790ghJA2GMYuRk7479aLYnjVjn8y1h9Ir
9yc/P6eMPo5kPy4l4WDqyEaUkIcyYEQD1BvVGAz8Gwow+ogF7hgjr0f7i1kOF7oHRyF/kNXM0f2Z
eWO294JwcvH32cJbxtIzqNFPOwpqDXF3DGjJBYM1H2kFymLjUMJjbXQAibWVYpJB0fhn+cikGE/k
fG51YAC4nWOHVY+4y44CghNKR5+stbpJ1WWl0j4VPsSzbUHU12auxQMXcWUjgTsp5CCcmN80b7Bs
hO6o2W31SmMjQu7YmTo9l8MR4Lysff5DZCnpZlBhgHebwJSI5LDj5k+g7ummaFx49V213NFTMaz5
C8aDRjZuBmm3ZcYlcqWUmeCtCfwmK2T/npB07ggVo1EW8twcPABnGXaHadjFIJCmdlBgbkLIjFjf
FTcx2Jjg2QTr89Oy8+NS6adsfgH0vtXQe5nNnGZEBLDZAX3ljfPwGXXQNY7E5qz6OBIncJ/L+Wj3
A4RbHxHVPQ3uWYXHDSGjBO9/Ukbz/yyKpuC0pkvXR1Uw9jxI/mAUWg991CN8sS9gFDetWUedjrt1
AIecIyI1p+R179SdR1qq04G47KNkaEm8Rgju05Vko4zebz2bRz8pfOBSdToxP/OvbNPCabTRlSxs
iAXElpe9v1VPgEcdh+JgzCuSWQdx9Uesyb2l6rXRRhslmBn/PXSpD1x2B6r8BuONFjO9ZJNJtReZ
q08Apojd2V2M03rhTnRCWTI69aBtUioZQJfiGe5+2XHS0WIexi4ujO7FihKBwNQvrINmMOFHtHjr
wnC2NF8rZePY6kl74mxMaXFAfr7U9g7To7C5Q54wxsku73JjzPWyiqdIDMMQ15IywWnh0aX2pjDJ
z+ilhr2BYRQZrGwcCfaa4UvgxY87TqWccYd45tgXp2LEBRL0sI6s4fO5i1cA05LThA5FKuz9Pt4X
RafsKBMgCnt232SHU7Q3PaNmA0aaTSv1CxgsdUNvhn9wFCMqIIIGruYPT68HD6Pwros8prJBLv8X
ZwxOqo7ixsmhreyIU09F15mhmZR1x+ebrFNzkZkBZr0jcUHo5sDWEKP6CAciXClschhse9MhP7zz
35Mt4LTXuvwqD/h0DoilWqX9HYbmApHZ/FHKDrlHKgPLSxj9n8V8v0YXS3xmzlg7ixD/Onm2usxy
p85H8mVFuIfu0dLBtK0mrE4xr6cQGtIdFmdZxbLBJscQCnHDerK3WUxwRX1luX92JEyA5B6h74I6
TF/KFsm18+PieoRhb2UviMSs8iAI8T6FzoJjtdkShYvfUqK5Fc8+oNDMEYsTHa9ZZMjfd6KwmLtS
XDQIbEWkp6y5bmUEdGtyLm66OI6SHvHuRReuFUq7i+y2a9V6f3SyQ5oBwFiakTrfbmczyFtXuu1L
6rBXVA+t07AWDqBEfdqNBO1rFJyZMKk7nWra5RGcXRK4heSW+D05qyrPGNgtHWnrLmWB6q5GtmcJ
QXUphaup6XXhoezTEYW58MChZtRd5lKn8QOHCm+5ayjhvlI69bF0lrrOoiFzpc8h90g9pHHzEHJa
hFMmQ38amG+eiPhd6YjkRP/f4r/DRDn2j7qrjId/kj72R53pM8xwPbuSDVnjtyawN2ZFvIgbyMhS
us1NYCaFeWNs85n5hS1IG3SRjr9PL9EL+smjwE2Y9N4hA/cq2A7EvxArIPN9E4Sf3S9Z2aGEbc36
Aono71tOpHvjTswZpo5r4ZVufD211L9yY6mXRC9Ve7d6iSPV3dfk5KsP237mkkJYDAvrpwrtfWjR
FoAdsx47UCYwRCQiDthiRa3m0RY2yw5dO9pHSY41yBe1diDQQkXkLLsm6ReCJTeAH+MPL+rFQMBo
8fKBm9OZvQG5XWVgLSU6WZhXsK38NZhSEWIgoPMchnX9gFepWRdbIkMoWqzUW/xm8/LMoNmUJuhj
s9zDph0lpwVcfJwoUpBoanJ3jjtpU3UesVAAYA1zJ5M7XPrLSLZC8KXSrASrn+5CjvNgVmbI6S3W
kCl21DNV/ooqmnb8tslmGsrFlUpti1DQsN9M657Kh+mp5nh3u88QNUSFrL6bAKLZr3Rvj9IYtutq
cN7pGSeb/FmE6VAgNCEN3+JFjMYue2YxDQbOJMNpOWnYIcUQnEyO/1qP/ryRiVkyZpdXSB2D/wdw
YsgC7nnoEs54oB39uArbuRzbhgUhznWV12ieteOO4IvFZKkteRZ0EoExnNgWpdQYcDJknBNndRnK
8t22zQPE5Ue7HMNKgw7LDfnvjGD1SPhkyBrpz38AULXExD9iAqJD3PQXoSfyCZVrj3SbcqD+yHam
GQQldqU1E/SmAFVjiMVWugis9tKZSCDmQH/StSsifDUlPnBOF7aS6m5wHNsyqbo3bpfm6dd8Sdlh
+wGK8xmvgwND6UKcBe5kgGWZcb1W4lv86kc8FzIphFPQV/tLGNMWUSpYG7Ioz/yCYzx04NRAfQ0g
fgHiMQGrj2hz6XfDDnQaSkAXMtBpUNdMdAfisGRhgdrZkz2Efl+utIHifW7XlokXBmR//1Imt8pw
Re1O9gy7udCZ4ISkBARqX8tIXywL3SK93l3IvQ728K3mQJwGCtksUGpkHoKO+lcp/4tZwr+JferX
GyFUANQGzQ/9reg9LmvMDGbLiMJVwLEJw4neKh+LWMLcYLCsLMfv1/IHWKHG7bJZ2NdQ2KTsnxkV
qt9cdYadWRw/CWA6Ys3BxvUw6sLUHMcjeWDBMeVlCJaNk0GYwDYzDKbCZP2O9DHTvTYG1NLONwzg
WxT0fiXibeAVxfRoNo+dIyJ4b1UCmhdwl37Mg/pxGchOZeAD2/lp7R3TK5rBTbTxE14sVgtggPL+
+svcQ67w6sjL0Q1rB9PXDFy1aDOcM2ThERHCU1RpegXP6JO91GRG/lyG5sRGBPeeMqlCJbC+7hbX
VGBrnw5TDBJZM9Pjqu3s5xJThzV+4VVDolNO1rp0azak9udVkVlBFi7akhegfdKpCGyIAJ0IWyNa
qYh2mx5V2UTimJnamCRyz74AbgmFORr/ADGWZe+hmWTxTiDHu+EuN4MXXT3abz15klM/otgFcH8y
Zsc7CamfXAzGcrV7mxWQtzc9w/d6wGQKyIPKCrGQmTF10r9gCBPg2f1u+OwX5NG1+XkF8OT/cKTX
LkYi5m6CPAJ+Ue4z1QRwsNwyA4o8jcvaQjOmhMxUgA0XmroF+JFnlf4ZPhp0mCfKhFxGXXHBMuwH
JY+R1obT1RPOmG+6cPuX2R1moBPBgH6BntbBaeagqtZW/ZMHvE217WRrdqkj+F4wJ59eBxFoLmnJ
4NlYkS4umXivcx4W9hVgBch2/vqNRgPnxGx3OCRB5s+k5gi/86RoAl0hGVXvVKKVnuHb1D7Fan/y
68xfmbBELKft2122LHTfJXbTOw+t/+mFdCOsTsA5jj8+Zexbrmp0h18svtwUcmHzy0SBHEuUUsfd
QwBaMTHaqz9hFVuvWFgU8Uh6pRI73PcZXP312wo5pJZHOij8wsnGJl9CuDg6PL1k8q6b1JDI4zgG
w00gMwGzv8pyVn75aFyBxDSCN3s3HLQjQJPu1qSzHwksdWHqn/x8RKpjxG15/UbMP/0Jlt/dwkJW
y7zZLZLEYZQGId/UYtu4eAkg9B8KM6STtgkKy30vIPw+Z4HfcCng6B8/hvH8zlO8FGrUjbXd2HMD
iRM0pUF99awRSQUH30YiA3X7at/5V0dPbj6p+R6sTiylYiW3Uff8F0h6Zs0vyzV7NEdPuS89eNLd
9smGr73jty24jWYgJpDzHvdDsDQEu5L02dgLYIXMxhnPo24zwCTuTca9+Xc4qW2TkkAR1QvyXvJq
Ng8IL5v41aQDJqs0UbHSMe3TVB7+/X4TEPtV/T/XT3jMD0dWvKLbHTV4djsYuwW+xcRfFaid4O82
X5ntEP90vCQkIT+LqDCdt5OlnyArkVKXzVP+JjZVROV+OiT537ftIylot9VtShmZGVvMN4eGDTOl
daKyf69zyqT/gmiTlH1b76+5okCRZWwQvlgiLgiktD0Os1EYwmcfi0PftIdChwXptn3aV/5GaEWt
gbGbHDRJ0khQJQikMs4zDvr94yaCBHsX5aXIsG5hJQyMD+1H0CX88rrUK00gq4DyvZY+Xi7Flfg9
zEqdXVuiaY5+5qZ9IrVGfYvvTdHgZN2v0PdWxi0Wmk/ZXH1+AtULvZJ8a4LqKm7Ep7tJb48jru9w
WmUu3PrxAoXR/6qnEH+geSNgYyoe5HFviyioKxc04hJ9sZ8UvgVbSSK1m2FWzDbscR2cJUdcV5I+
U7FiDFGTPJWnO63hAk358hTU0gIo7Nm7BI85aIQQyxiM3dpuZxhRBW5CqQNbIbA8hKWHyk0vGw1M
NYeBasoBQ1JfXwWgolRMY8gSlLXkh5VkvkFi5S+ZfkKxuozhYt5hsJ3lLTGby5t1dfsQXQdDnaAp
6Q6z3urktgZ7KdpBu6o0ZvfvlwCBamtPR9fN9hQDCnyqk4fVafv/f/J8t7oNUhYU/mukzCQPQXn+
c1Vwu9EmkcBbNs+zMfzJr0dGBqCCgajUOAUb1gtVg2lV+MnyAFcDm1V1BkqK8ofPkDPRTBeShdSs
7sd8SIZ3eQZ00edqpCsB1c8RC5mp46qH5RJMnzdFMCBijRkV64AkInZ/R3Fv4JObRbAjbV3YPcRb
G+Ra9MOxAJ/JGy58FiVN4qmyBo4wCW9srtj8u92NT+3iBehQv8CEsR9DFW0gg6H7nLMpkB41OcZx
f6iBEL4KYFUpsbWcXTfdFc28Tg8hxN65UMgLIybIgzXQPL9+NIewM2OS4cnJcn4Zs9TGsDrY2alo
YY2vTPsqqks9SpVS9+4ldn+bOy05C3hKVfjIBnDm72xt3SEFq4KHvv9F+s4K6Emtv2oBwANSZEGV
E4ZzwqeC1NyqwGgGvp7Ol8E4F9Y6O7UYrq939HbLkPvPVDNrQS5SJuDbQJlaG5ve3Ol6FGPGh6km
NtaZhzJJtq2ctiSfDO5bBSXGnkXF3pfD91t9NZk8wMI7jPpyQ2MfhsL8vNXg6rGcfZGuTs/ensVS
LCsUxPTkJa6YtIGq3bBJr2mwSdTRIFPaOQw5S833kXeBLk+DT8mRMNvvlavtDEPhvWc0ENNIbzeg
zlAo57RwmmF/4rC3y/R6qHcxD5bYZiZn6myLo0kFiSmRSqZwK0KXl6mOfHypfuDp3GLM5PD5szoy
8urMM+3I289bGQlrpWucjVMWSlrEkdqkSv4DtXnVKLHgKa8yOF7Tjje0UaoT9AVvusHCKY0S/yhV
OtsdPp/pJ3MBnNNF1Ev4QqkgpJdWF3Drr0+TpPmGU3mYxWnWV2tEDX+CCuigPCuC6MeOudkzmWnI
tTNq2p/OeDs/MpdRtIbxw4YLil/tn+ilq1svx9NPQKEFDq76w9iMdDv/RHvGLjKhN6NdKLIrjQIl
7ceoaUvKMvBTTKEYmbluhlnQOKdmE1qzqPXDkSET5Fd0QNyubazuaLrSvhslZu8AqCsp8wDT4iR6
baX3xVpYAH+IXGRS8cz4CkH2SQ+GkgrrViG1DwpGwSMvjfiXMxNRkybErTLBTvERFLxhopKJbZ1G
tXjCCBMAwKbKrZd2FfkTCK0CrFkrQcPPUc6QP6GXH3u7DoV53IqlW/74NA8LnCICx4ag65yR6vr3
wvpYnXHJskRywZ+Up00AooMRtPwuqSJN0JpHa6BoVyBNjCqKciyvRP2SYKkeNTd9NpBJtbmaawyP
ZnnE2XRSXLtfTlNkbUMbJ8CbFGRoQ1IPEZgqp8fP/1uEvY0a0NE9TTq7TcdJl51511UMZPaolxEF
A6GzBfT6pOPrnBkJyUWGCSUO7L5nYX4t330ZXrJWlZoPQKp6A6zkicQkVIrOVsSVi8jTQvWo7l0Q
uvHTj91oPCW90ygZ3IXejxnIUI/1abPTOvivWztjdqU1J2sauyilm2AvWfOTygCKA3eUomf5tVL2
Ohf9ccrqIYSns3f2QzdFX9OGE/POB+SUJc6ob1r4Occlz+BbfR6aThq79yHSs2wYZImkpUdhFCxU
DVjbkpp6qvbFxzsP7Kbc3MEYlLZCl6AzS9TbDsqVZGkcuzgTObskk/JQvRqvuG5lSE3nLQ2kEhv5
HUHlYLAFJSG4Kbc7TebWKr6id2Xh0uHe73mcP/wEV4GBL+No3ngpg+uHpJx/nkUTLKlphBgTkG55
1a33Fq9bNbhVME/sBrWfKfrwVG6Op6fMjKrd03hzbjQ2hLq1p4D0af9k5xceuoH6BArWQ13H57kd
P1ZWKNvkEpfbGsS6MuzRkOK1A8SIxaDr/ePFXzmRvntxn49m8sqrM1dRe4hbuJgMqDV4eGt9uPwl
yULcbzuLtswX3l2kfuymsJHlbXeGfeedJP7eNzYrb5dRWMlk5VGwpd8UhyOL4h/WCbs5ByPsV3WV
5Ny+KPPPAZ3fwupXT8PFEClmb2Y/RGHI/9LTbleu6cJ7/7HSI/Xzft/E6Cvuze4XQRT2a5Dsg83R
BrXOdq2ugjIS3qZzPP+xzncgGOaDngc2Ckl9EMwm0GWaUlnLR/9VcEu1g6esc9NUQ9NJeQqV0yWo
tKeOEThZNJBtN7Sn9NPKNxSNX+1ijF/COiGAiSEdsJ/aLBm+nuCHCCp2q4pzSfoyxInadtp9ET+y
ZCzmISrwwCN4DleJdhQYs+M1rzKo13p6AdBOBbXeyG0rf2qtIcCKcthCTC3en1PlvIFpYWe8ijf3
yV5loMK6eYhCMfmyFUUEEJWUROdHD+TZeUMxUdHRQSHYSTKII9GD5zXiTHkuC+R7fWuOBMFckY7U
HXIEXQxwTnA5IriK6yH83ErEeQ1CO6kG1k7Dm4EpCbh7tM262i88vI/z0TCF7hp2BmTWVbdg9rbN
1SZDk5v3l0gMQBz0NXOey+ZmKEvSYVOav+qKQGzJkdRRd2EtUWzqhFOSf0uwzy9YWpWgnpzm46cy
6n5j6QKzDi4cHxbkfFOc+QUUrVXyTaUCAOjHrtg/MqfuH6ghd9SwkTBIQIzvP6z0GUNUcpd1sFFC
l0O2JhqU+lrn6x5cG0sg3foSXDhOEnuree+Xpb6hc7k1B8Wo7lpzUN+7Pd5AQm/AbnacMThRwywq
FAHNvmnYpALtnqZ6agZP1YQeTImQGcfAjJBLvYogJ3nPTp7YMc9EkZdefedYdP2bQPgMUFgM9F6U
EfddA6WsAji3eyrqW1yVCFmu5XAmSiyAJKyIdA9U1wgrg4S+hL6QwYD/92OETZG7dow43KJi2GdN
Q4mWxWqE2VqNuG72jIko+H9E/Sx7P8+RKgLFm4lJB8hkcPeyMggPicPfSeBfQOVYjYI86ZGV8eIw
+k5SLue03gnfsnzIRwac2uWtiK8c5DvnbfBHxGZMFcMPR3IThUktux14l+RsSMMCIDO8QDqm8NVe
jyYefz/t4qRDQ/8ES8jpGm/nyhpUVFT5WJLwbj4qnGowpbCwaV+O+euM4zErZoBNcXFYV2X1jvIS
ahGWpGHSIlovCFQM8DyS5ogB5uygdcGamqgeQyymDs1Nv/HdTFQTbmC8B9dO+HYuzzm0V+m/eDhK
45Vno9ArQNLu+ihkV1++9CdcS3gCB6335TFQFPDZKq18v7DaaJHy4LycV6C6R5yMANKh7lb2KT04
K+eUXL2zo7B/vxH4qpx241A7P1edCN3bs3htwMpluUXBrPmXN6/bkhhGuK5bWJQ87vDQ2xSACFjH
kBR0kZwGJk68PwyZbhqA+gY6jCKAtZD3DKr0neobzyQ8DoZjiRxX+gN98mAmsSIZcHvihpqkNHPT
say87NbZScUKw6FpfRl23UuQsF3DfOVicfuG1kWL00fPuDAfAII5us4h1YUEEXAIbZTH34U/yAU+
Id4Ld+voIhIQQVQ1fHgROtLrtlYoVxt2Pjxxb5vdIi8Vo+KfRr8RdsmH+1ME7j59bdMmY6J8XELa
B9zpYVlVmnpKRM2zwp9ABHUL8SR/W87ZgTSuzovQCKKLx9ssHOGDCZkyCh0wTHjKEBdWKITCboum
af7caMcYIHx/ZVy+uafuBjWgiH3H1MnbWnN4YMlzExzfqQSM19Mgj34p66l+6I/3z0BPIZ0XW5QV
ai1q16eZLvLjB5oLcTFt0FfRl4XLSgWD3EZ4jlNwfA6lM7Udp/sF4z+9M8Lp0KY4qMnKEkpfxq+D
1FNi9ZuJcfNKzEFRF+XyZVJT2EMjfxe1VKnEX0RibSM5QTx/zfKDeYpPjdsCvdAS4OD8ULKMdNxO
mZJdMe0N947qx1iIfoBopQmlp2mRM3JBWe4JojwGtEgRd9vP1tRpzkDLsCzXoxMlj0pw2JrDMMe5
fdibhH7t0531O0uzLnA6vYg9LZlEZhFJg1feHwtz+kj/Q0mIX/JNLf7JRLh2dBlIJ30tHShZ8Ymc
LTfPBBLri9jjYA1UFQdFQTLuMFR+Tf74g+Z0ya6fzX3QXRc05+XCYmMkKhfv9Vti93JMbmCfJuEr
/epgT5FmQ7GiqpVnM7ixcM/NY4NskadqbEUydIjJ6cE98U+3nF0Kz/cj4UxZcvgVVcGMmf+ukz7k
rTB2EqVktlcCnGeP9CkyQjF5+/fh92cRirxVh1YIaSIU/gZ/YkoDMMlzy7Of7/2mC9i0xLVaK9Wh
f6G/Oj6dgC3duIATfxSCqb0LpYCwADhL8G2o1/3zhEwlTMdDvInaKDL8ltcY2dSKjOO6Nh7n7n6N
ZfdgVagVdMtbvTjJFYKcr1vEHotDbouHtvPphwakc2Gk8eSx8IyBlBME5Xn+b8/h1ly3P0klhvVZ
R4Nc2No9GGcZC5nmA1408KFSGLRLbqCbSoIBqFcG+UTS2XbXk2HwWzgTw3abCIESXQhbL1OufqGm
6DFv1QxH2NWdFMD/+P1y/JNDnAr8FkiNpifSr5LkoS4aeBpngUlaLB1S/X9n9JD+O3at7+k6dL4T
pONTO+v3YK29pS8j2oh0Ss7KB+0yzmn7bhsKGSLR0VeeNKpL/IjD6FknhytcZ5SVyf0Mi2Y2A3ev
S09R6fXkEJKPP8tP6hp7vzPbZGBCcTs3K5ukE0Lr0xGlhW0ssVx6428dIv4pVomCCxN4EcWISsZh
rjgvuDaXi0R+ki5KawU/ByxzS+4hAR+0IIPu2Y7dh604tEgOW44Sj8oGPzoRmT8TGXAoLuaBeNDp
77RzYKVaG131e2z4s/ZvjuDndneSrYABBscz6p0J3Zo3pcFNoaTmJFY8QGAN+93/CZUoriYTUJ9u
cbBGhfFUTLvQ/MPS6wrK98kQB7Uj54IU6BRO4+J2sIyBREOzNSy/Qr52hv4LOKiMz9zyGbExJwB/
dhl+ZJUaIav96Z6812yZUODTlPABBvLaeutIjDx1xZIc1qOHtIkm1i5Wc9J/+YsTbyI0EQ4Q8OCL
MNYAl8PMq++FZ8NQYcxv/sm2Iu7/wZxk0z1TSwgKLowVbRRcaFu25a/cQSHKYrrY/zQodPItdQAX
/IABjqSaFdSmA7pHm3EcvpQkHwr5rmx8cTrA5cfwWaRkQ78i2MdAwPXCn9WE5W/1QQW7lOLvwbJu
A+KckcDHIX2YvdT/AWBGUUtt3H/UIRvpY/7dYxBzYLFkf7t+QSDCh1VeJDfMrCuYmC9DrZ5IfBsi
F+8HQUz1TJ88EOOMdB22Edfjc9xmQW+Zx2MEfBvHyNorZGfyFWeYc19G+iZLHflIcCD4zXQwjNky
kvm8yoYXDgXp4Ouy+NgF/ZLcNqxORuoQPHqOk5fuhIVyQXix+fLSd+QT2YlMYhcw3W5r5jhdDfAG
z2tUVXm/R45zYX+pCkjvk1JbLbKcVsz2B/dPjeFQnMvnJqtJRFFWmd6NZ67Y5A847YCHW2JegiSh
AU2J9ZH7A9Cs/pCgDPjShnCsw5bo8kWpbIh3QPU113c1yHtcbemPeyaxns18CcwAnkgGvnUIB7V2
dDNuTECX55oPk3BxZmkWSAk2Xtd8fnabuTxiyp2dCArFM9IywpE3l8MsM4/M9xyEj1qnhYWvhpn2
m5do0+0qrkH/2jOhtlw/BUJfc56KE/N1X2YRWiuWF2L2X1ph7zbl50le0pg+Zer3PWpBs42NNm0+
p13ZzzGIfiNyaJhnamtqznXjl4LJWFT0FtMii5WwP14jw9LSkCbav8YFL2TNzdhgUhyrmIGQcd3+
LsZlZvojrgw3b9P1Nbmhov+TEp5oplzoafvNqT/isYqUZvFLWVFbMngFG5gSnf2QxPIrR/R8ndWB
7s85nJai06VXpk6EGogy6sgml5o45DPH0tsH5WXL++ZhejZhNLnOJ6t9Bbw94CKwLyq97UKw6oLo
mxMk2VP8mJwUZHPflfzRDwyIiqkpQKvfGlkmYbpICHb9xiWcNM6ky6rDRVPEJKd17agIdLDLXpvE
h2bzPbmXKFX0c37DZwcFsvhEtGjrxrTijjRrSPRdC/uU2Ww3h6C9WhzQsiE6GEl4PaiD0hLC/VN0
XlG/IOxu1c8Occ7FdCBbnv4n9XUnNLPFMvoWVTSPKS5RY1CU8+heMJViAFU9kskxsd8xUD6XEM//
aycFWWLLVg/Pc4ojEvcbcerBUdSPxWPKSB3WbBfE2SG5qzjX0yDl+QFzlJS/ulT4TXSOL/8KLfnC
ea+KNtw34b43CN1Etcs87XZTzDMe6GS0+KKLOqvK9IOabIU3x+/Q1V2jMl9PgHqV+Ahybmuh39y+
8lk0YNmW57MNjS+zjtRFxN7PsYgVGBzbvFijuwYuWDtzg0IoS5lTMDsTtVsi9D2Nhc8rCNVMolrs
SDVD0NedhEjhmujxjR6/4/yz5y3H6YAR6yVewXcbCq4CpRcdPlP1BLHCN2Kea4MFlnNApm1TQUAv
IUXUwtaCo6bxmVYnemqZwJu+VDHdRaYgSJjgReC7yqDZ5InH+CKWYz6MyckQcrvCBUFQXZEbU1Fk
8tZt6qm6ruOTrcIp8c96oV3s8jyl04IrF9S6O5yPVBxre9BTnM3w+2W9RYEbJuxNV1m9jGb2cCHl
XpKUCC/XuclVAiV51VNR4m0EFXv0ghaSr9eOTUOn4a7OVKlYkzl5z7pzZG13T3wh9SSJIdQ6soEC
Z83cO7bisWlOj+HyJlrcXV8qrJaA5NwlFIh+laKb1+CPjS7aZwyZCw4cGBZogpVgDwqlTVDet3Ul
iBIiKqR4j57Rmfk5BE5USNuLbTqOYuUbwIuo0fwNHxat3S379Id4ax650zIblA+GABdA/lDQV4Qj
WJnNPrMWA+ObraY24VT6J9boDkm6vg1XjDTBkqx89Cow1oh0QS+eIxawOrOF7P8HS4kMQfQ3SVno
pjCzQETpCr1iIr50hOY/u2FMcUL0CGF8LKA1fJ7GLOAXd9ckUcdda/YzMYzOvqmYaVuX4iURfUzu
vPCxb5TDcAdcXe2JYRiaWWFrqm0GaYmMDZXc/37S1M4DDY8lLk2SQFSvo419sYev01ZTbz1lChWb
7ORDXPRog7FC3aXZ/TQlpB0J1332bnFMF398+XfeEqhSegFWTXK6AZ1pWzuHwGjtif86mAFMTOR8
RT3irWSw7N5EaPwCn5A3cTGvilLVKbix8nvg0tQNrB1HUSrfzPd+OpOW101FcSNQ6qh6Md+cWO6C
+yC8yX3xocC61ZN1HHpCL6m5AwW72ZZOeI33HRdzw0hS2akAF7cT8F9WIkkZVyt+UvPTqaRhVawK
GmjGGo29mglxxgIxaTVy0jtYYhXZD64pmmerN2p6KqUpF7UL6W91tu3HV1afk1J/toE4TDmAddKW
4EFVWMd09qZz6Td0ATnbotReC3ojJgOvl86Gu9+OonTbyGlUfb/t4iDDCHm7jcpR/QvcQe8s505m
ZfV1FknRkwPf4Gg6Du8GKWxV3tYikXzJErA1JfgHMrIFotwMzYpWnGlaAojWDLU8HZiHPyvQIcsZ
ed7/Atxqq8jmhbqM/emwMjbZFPU9yf8BC+TZoYIvvVwKuOs9D+9UqKmgqNsOq/4g5URRdPsF5Q1x
ls0TLLxaY2+rz3zrS4R5rII2XN4ND8C75sDrhsm6gK3HaUCK5nLYmmpbV1FtIcLk3n9NrVfsccIL
MSIpS4imrbAwDPG50+/SAjazHfmLisaq6v3e/99U14zac/Oxxe1GbAZCmQoU7u3Zi7W5JpCyOhZw
z/QAzLqXtXrPb4yaTsaZnu/Yt5suicRWVGQtaqHkI62RmxwPunNJBvfmK5B1Ia8sdYyTSkEGvG7b
s1dYilN1gUhVXDBQjspFQj6hCjFzXyKlITDWINs+1GPfvgRdyw20cm8eygJsu3s4jrt21Ytf9V6f
+gfWTFRs+qUo9iUdFsmK3x9J4t/VdMuesZ5KT1YtF+wouZtSM17tTBbj8wE06sCf789RlRPSsDxr
p1iabeN/zo+G84Qb7HHskzBHTLRYAPu37Xj57pSC88a/rMI0HaSHGeUpW1vioMl6E06Id5TOxnYl
qzZPv+G7StDJJglpDmWasZ+uCepFSc/QTJ53lUEkrGLqBFDq76HwckS/9RMXLECQM3B0IeF5MHP+
tCLEFLj8BI9pxJK1rFz6Dn6RUB1sP3RsldbmbWXah95UZc7sA+kGkXIhhUXxRhZ31fPD+uZeKdn5
HJ3tAwiHeTJ5LwmcqItnuxwU9lfVG5uSaZXhW1uFijTmPz11v2q9E43bFwiem44Va4my19F0h29y
m4N1zzkBrJILEs5smmaqVZesJ1C2yEgCHGIEvcsxBos6GGY8bpPZxxbXHvisUK8f7q284PdyMclT
MhmFdZkYH3o8i2JJTZFaENtBPj9fybK5AqkcVThOmY5LWi/BrMWXzHXCboTpIhzK1SxvektOerHr
UXAT0o3g5bJU4RxmfBiBmCs8IOggugrcFcJ81i0BCvToZZt1EAgemPsR5ryzly6wNI3IfceNQMSb
xTrbHo9LfJ45cq7hGx7XN5bqPVX2JLfr/uGR/toHxA9ltoonzb1BVOdcKpIrDl2LmnT1B6p7Mp4z
J/A6KT5T1Y7htdaigmzk1n+9GZ/73t7eSq4VDkm2Yj9RAa5f/Y/d3slshOgb0jAmR1TU6YW1H26M
uKqOB8aHZ1PsFDJfrrmrgUJ6uiacOpxY69RrI6GJXzr6k/vAQZp+Y7+Vt2jyBrK0Oni3NLso0eQP
6K10J9Q8mv11R/fCJMq/RG6xnfM896aoaiaC0O4FG9yRoF7x1zpfVisTNE91vQNnDQWAsgahe4Gv
WIv+D+PgyRcTRYIACK3PuAXo8nJCTziSOUW+/lX9TnSdN/xNjm+DKmk5XSje3O79W/lBogNjB/BI
+w3i/Dxtwa9WQlTIcVtI6jfIQH0jp3Nbzj18a4LEDPu9i4g2d1fZc1m3yxpkKCocBXWBM/3ynVJv
T+1oDmMUPCsijjnYhWhe8u3U7D+hBgZYzQTVs7mHQ+801Bqc/Xnjklp6VuDs0/MJJHrg4oOkaZZx
lMgci/vDVt2FcyxVDgN2ehtIi1GvoIn2oec/f/iwKupFeCHGMTwS8LJ/v2ES9gViydJy61eFxllO
3pW8/spfwB6E91bkn/naP8hDsYoKz5pfg/ezoBU8Wc8qHrNF1EfWXbA5m9a/k7bERo8yeUPlvgEw
AqDQX9TMKwjr7Rc7nrPcumXa38FdtEioqlWhJCVbfM6vy4h5y7cZBtxNAfM6AvGDs9PxVD+p7BJb
o9SyMn/DrsQnWP64u/qIYF/3RA4UoimhyGhR8bBdYg938FcW+99Dc7EClaAjEQ5zV4xk8IbObmt6
JEQ46rzUlGcsok0VFXjfFJAWzbN4l3NImzV8I1TTylJruBXr3qBnL9CsqO1FABmGqVucA98+Scw9
2rGZJDOBSjKDJrDeaLzQa1eeb8ekaKCNDpqIm9LLyqCuge210kr/Mm2stPhhHLG3x3GxdkX6JHLe
zuWSxNTZhVC4Cd9mvm0IxZUMZqzeO0RTNLz2TJGkqjEYdlrasfCVP2i5PpNS0SdZcheagoxpk/G6
297ogRsC3lXBEz2IgcWVnb+tnymKbiW7BayzipMYFYFNdY/EYLxrKeBZeHcBbNltfWrt5ESFFADW
zKrx57sXJRrAWOIVQ8NZqy8V6P7bzmCsObsTt506eNEdO9F9ftkStz1qhA+S1VzqFc6vReOQVeu0
rO9e57DFdRc1kqAmjY4TbD2l3BLAax28zjf/OG9K+2mNvq0gmmlclackt7YW7YDVBLG8NFw+gACT
bQvApp9zMIxdMNiZLHSn5aXniV4HzX2w5T9yFm4lBQ61Uq3hgfYH+pqsiVbeMkVkb9MZFVEOcbU+
g8Z5JRDSWn5wtREM9XoykKpAZ2IX5z1h0h2j2hnCAWz5T6UVdLXVnH1MZg6TLyt/z8+WbIDNc8bP
UZ8uAWkZItGvrM+Hdbs2mXQSYJxzdsLOnq8XXh9f39GhKjsjMEHE5DAkPBh/Pep8DZbDOvoj2yLv
FAHtsHF+m9oC897OWFSZEiW0ZuuMCoV4lUKgvE4ZNqgPvdDMY2FZM/LEONMRk8jeBd0+UW7hhOit
8GOaKdm291SLt+7gm3Hrt62U2SyWkDhAywcUTRpCQASXAfEgAD3vd2gg5b3bzjeo1voW9IPC4gHA
070CnbpnDjwn9BiGJ4/2vjGnYHGlGG/zE46f2/+gfv2pLBds2BO6EUrNsrr41X4zuIW7rben7Uo8
/zxqRZn3rRvC7cYzO4SmsJRj7zgUt7xAA7qZ523gj5PZrMvXRlsV9lnCV6y1m7vRMK7JE/+T/Mwx
/NIVhgecjnJZG5MUhsUhnhGQ3OFCWSzR3now0fNb4eq5Tc72wfsuzY9BqdrQUb1w1XtSNAbwvJo2
lMeySkvJuLN0It0w1Ccw+cF9jfyV4ypowgBRhYCgCeQmwAMaXjR5KCWFRPbovGqzvdgnz8qdzK5L
kgb+LInOPQqWEC3vejj7EA2Ox22MfOuLve5EtAvmyETr+xFFWjKGWo6qZSUgCIqg/XQ3NiECqs10
m5q0p6vx/IFL+WHYvLuZKMRPN3EOny9uDUpJ94x+y0RvJB6liZq5aaQxMm6l2JDYM6dqNcubH6ie
MEDn42ppUzgUNJbhQQiBWfcSp0CzV+m8eAHZV2s+U5MwgyBUeSE2pexWgrAt3RoDs8aU7MTLihdr
M67eyAEr4uo/cbIWxMV3ogtkwBroKeIB4J3I5DCPrgbBTGreiyljzKV/dhuyWMnbylFmhJWS87yT
xybTRo2fIcEYS49qx4tAbFkfPvH4tB8b/kIo60j6gnoyfU6d3Z+zSRNGo3rsrvT9wYhwm/7048po
Xwa1wcbYOKgsgF0OhiqURCHpaZahCfL/y9j111XEdFn2NEzKwzcgXyyav6MQxXG2/CLPbey35FSO
sc6BPpZNvGiPJOW5w58VcK8GOmHrySl7PfHyKXTiMNTvOOgs9vkASdudjOUmU/ENCjKVeXSgax1Z
a+NuxijqdOlwdQVmjtYJd8iH4RiTjadjviUEsLhuUA20JUxXVhrYkdmEZdmWtxKlJbEI4fGtco8f
VFfTTP4dlGopKP6WXbKcgj0Q7hyzscfV+Z33+49EX4UqsRXH5kf2vx1BqMmy7jYt/glyMLv0f+JJ
eoI8dNq0mJfZYqzhdw/jjuEXSUgN3Z+56SkH4yPHyy5JOsxSJXGBVWj3SFw0Kch1F0J73b71b4Tm
jR2OBFBksHyIDh4HMH/piJRwsd0i93kClVtbJ8gzPvQ4Y64rYMqP0Z2QCXkPydosE7Y1ePuDG+l/
WwbIAZB4TPbh2KtqI6PNmBCj+1I+eLi2CTWHCFVnNSk5qzDbPF88788jp7GeIADlYI8/aQmJhEKm
4VpN+yrEEb7/fu+QlYgtnKkIdD3avaT+8HsUhusIPcuQupeWxlFHf0YctkAXosvdZRK4hpuK8mJv
e941KB+tPnRaiE0DAO7oUy/OPGEwVUHwyu/IbshTCua/Eb34GLkvElVlbOaA9ZgtaJH4UJ3x8f9E
ARX/6svxt+BdCWrPaZAnJ2izDl6g1PDZbaH82q+zQAj4Dp2xWjejEu7MueW6SWy5qXgUN5rECjxQ
6Totqgxw3ycW6hLn4iX0bDW/LIOpspohCM92cL8AfGN32QFsyhr4jGyUfExG/6Gw5cdSGZ0HFmHa
lt88Fe1mDGMcNp/qv79h06bRP52NzCV53P7lVVE0KEvtwsa7LfWQAO4B0AbXu8Ikdx612U+zz2Sf
XpHO2/sUTI+jVvdyo+KmjHcrzqE7/W2nJYa7gaBwwIeP/x8BoRKlcqECcHoZbllQVTFtZTguLLBA
uhUBNAeUte7VwVbZvf1DoWxCIcPn9kcdzq3gfx8KL7xs2o+i4LRTHn1QUUuHb2vyVTxXFnHzTsk1
/FO5B0M+JP0N+ITkl4YtJ7nfx/+1UgqSLzTSPjip9LP2NgshwlMOfFfOpsIH0jUtfGi2LgFLQKLy
W8dpoa1bYuCdNz7Fc7uJgTRNKgQjScZ48qKMP4QjYN42iRggK2YtO5WaPzRDtz48oqtmWmONkxRM
R33FpBDihx6wB84I++QqJrlMFzKF4GwDD4Ll4fUcyw0BkIe97m8oLlo6xG7dkwb8cCEp3v0hHY2n
L1W/7Bi6hpoSPQTqRWKgPh9lew81O5+nuAO93wXcxdMwLEKtGJ1HOb5FUUfw/onoftW+9lEpDyMx
rMpjrBqe6ltTtvKQrz/4YP/CLFhwkcd7oPKavkXwrX/4fj2urvlRBOVV7FqUzGJ2ggbY5/M4kt1c
opzZFIQ1bm71MlVz8S8gxrDTEhZrrr80QGrEoTjs8moMdv9wAqi4j1Qwrxci4p2XLttByDXbJr7S
uzktpcjoQ7q2D8Q+crHPWxM6y1ogWlFhrcmD7ZiTbAV5sC2511dZAt7/0ssgP2NByLRyGNoQ2nNz
FVSxWquz8PE9V7m2BBZWONkykFVgBahBNXdu6ThLufWYwYjMEhMj+dYWMp6pVPFjdrIrdU3xdqkF
WcP/e7ToFQUfP+DWTEELa5dQ7zVaYM91FQh1lWDa2BN2z7IeFPXfFLsjeqlDJ5sPoZTy7++2hsGU
VyhLBufMnErEiEC2W4vc+T8sAsx+JaI5GbvhZPuMlhxMPyJyCqHlHJVajZ7SJZ8nz5PxUqNcsbAz
mZ+9Vb5tEus46AL8cZxJsfFw03G5deuceOAMrkFiG+vvn+GUKmoptMI5vie70tFK/FABNMFWNFh9
+vQ6zHstMiVoHUxNUbNx41WWCarWAl+4egcXoT14REVjMbpx5SoLDwaXzAOmlGTXYUrtlPwtf7WT
WIFSF8NaaBTv6YdSeyQnEDfrZlGtHKXA3f4vois/KIXQxtTG5MzwWLpGSLQ5TAaYqROYdfhHJO3h
VRiKR6zRn6bXqmnZETIlk4fNUxryHkv4xFvFMo/zEksxhChckJoyKZEtVsLVnbR2LLfqyNSqN8ZE
meh5d6UM9lEXBMVls95LBCwb6Na34Y37ArY2tWCpeY28lrpDB2WgiRsq9QXFHhvzy6QPxVBVhC9C
Q1gApYbByiFAPBndmNJrjERw4yq3RV+HR9660CIDhnMyFFn2ajEEDlKkkpFfUlwr67uuGOMMG5n1
XqKJDlenW3sL5XV5rcVVqvVe7bNVXfYmvNnu3jvUpqwVL7W5e6TGgE+psAZyXBed81zFRFicsUzI
LAt0+3cEYW5EvrTk9mSILyKsiQkjs/wgjA2IM1eT6sYDOVCO33kZAci3xk95CYTl4NY4uOR/wAWE
tVfKqrVEuQFrsCID6PVw8FBcAcLlCUuL6DJ0p0hTXLWcauRTjSFikItU/TtSN5f5HH1UvJoY41TG
vimDetuzib2hWUrQrJ5IFqNcDsibWQfsy/KQyJB9iuYwJMmpKg2Lb5HSog/5bjd9/JlMpkBWuBGS
adnQwTrHY8wp7E7VkKzRIW2Yk920hsMbRlvGtjZoV9LW69lKa8yimdEfdrHYnE94JFRMViCjEZWS
PCNgbnYen8cQj/UdOgFQ3Kt3Ykn2QFcqNTV0YCxICbcNLBqhreZvrtGGt45Ag/5O/qXp8Iz4NQ1/
qb3xp7hF0Sn/zfMBS5ux57wH/6KAAjQu4vgzAFHAbVOve/7jqGjFeBltomPLpJExwPqV2w+SZG9y
/vJ+3TpvNyELI7Bf5VlfDz4DV4wa42gGKgykPbiyh94n0Qrifha5j515ZaxaFB7nAl+2wbX2fACI
P3gvvmLz+vOAUba/K53K6v5mHqOLyyXa5kVRLFJb2MVIjf+HnpoOLshgVpMYGbgucUgjYIP65mSD
kQ5W6dvIduNOVBLBc66VfFM5zvF5kbp8QyvRhLb1A0mUHjKVAzuaqUdaffK1UtuUzE5Jh22VC4Uq
JcIiWHUS0t3YJNs9hx+S7iDpmIAw6ceroRDgpeo89g0rqelyT4PRM6/V6S4w6KER6jPAHOWVn9rG
tfrvMhiFXI2NoX9SP4Dz+NKRoZhJYKBY9t17Arl8mV1fOzgfSJlFrqjW57kW/1ijVST4bMasUCvd
qj5UOZodZLHuFMgKS0NLMtJFOmt9NSqaEWa6DrSapNIZ02tK9aV7X3AomaDgbTl6bkAhXsUKd/DD
RI8BEPZFGaCiCRTDpVA7ffZlEN3/fY63vzm8Tiwr6id6/Zq7ovrsSd92+6UUPF78nUteZNWKF+1t
HyBJ18ouhduImtAiWi6iO93yYsrGdouYN8Smt0YfxkDfszvqxry5bTmKi4/BeoZB+asyXga2cR5j
iOSvZbSfCS9+45MAYytOwxyXX6LhPsMxIG2K2O5F56/M8hAWKilF+KHFfo43HP5XV4gmaX2aAU5q
Qm+QeYXtk+c65wY0wtBM+uEsdd92pKRyJA9pbmXh0+CU09fQIae3oX3vtFdDfxacL0KjWAbgClY/
Rm/n5ucNnrZizgW1TVQzZT7AWUQPE+Vz0r69fgNLJLrDfYDWmjsL4eX3yEjWg6alDn/xjngMgwaN
XRS5jXa99ZYgHsZWOPk+3OTWhZs/dMPurx8PyJYxg45npSfx/qhnFKOQg0YICiiRjCLu6je40B2a
AydouLpsFfJA03TAHrEhD5+c3VCP6VqMPQ0D7a477lbPKsCIC5quSKlaAkDCo//Oym88+papSp5M
CxrPCl/TjmFlYG86BbwmLzmPOGTRQ4O288eRrAdVAswrPPfvosHBHcDe3kyeVQcOoeVkEjT/W3Sf
UitV+rXF0x3kfDudFZHyenESCXQ8opdMDev4LW3nYVzCEJ2P8Qecb0/XBazpynUrkKrLph9SgSsb
6tTETAIrK3PsSscMfqYqkoxRSJcYmRjg0poUkaBHSEKNSV37RDvfzTXQC6QQiakbuM7h8x0AKcQl
YXqm79CRM31TKQOn/ZtEMC2C1dVr25qxQjGvDbdlm80pta8RjNVVdiuZBE9ONn1h7ZOQ/sZTnTwQ
yFgwzdEjoJnVNgbTjCy5UvJHPw9W3XsXWaHvnkFP98lubxFVeq4UpC6rWITS4v1x6yAvafVKyP3X
/pFhIX/mMrphNxTmxiW5wfGtA9H1/ubylfK3LqzSXVlspPOxCNe64Gtt9NPfEOF/y/Al/z4XRF0C
0FiXqtiQfnlviCJhFz1RxEYN6YFDvbeVm5vEHLQ4lMzDZw/QSz8CMfcNsCF7N9c8LAdLsYoF1EdX
K5EtlR2POqf5YJ6XuVS2Rrgkf3LaaeR3EVEClhdsuNMBe6XPWJk+a4xZHuDS5KyCxBXA8VcvvYkn
GvN5Va4q3k1BLRiUwYYlYMsjkSUaDgl/orcZ0OVKfrWV5olBd4ypGxGzNCOwpqfOJ6WOOlup+dUv
M890EgEn7xyy6toktfrM71fI8nSKrEXLZje7ibEcefzRXiq4/CYCVc+PrW4z2LJx46crLzTGZFL7
0Ai9W8a2LTXCTFxRB8UTVmVY7JP6o0YAEzc2hDT5rZmhTEJyfhsDtYNjnQS9sXjW1NjEMrzN01J9
+il5zOMjnx9aE9Jc1EL8g496ru0pmU1dN7LqteCiIapVYtSJLCpLowcQYVYQvkHpJPu322QAMA8T
KsfelyXuPOsjkgDVWPoWHgbtncMbwAGjrJMSz2QxMQLJu4EyL4JfFamdubHNGcyrO+DTVp5LxS7S
+DjhYus+OnsuYejwRB5sjwuz3nQzvC7W4Gl8FplCz1YE4t2mvs7cqee227tdwqMw8qlWAJT4p4y1
8MTqEk3LDyqYSgpRlUfwaXzrneJAtsGIGiMzI82VSyYdo8rlF5v+t9IGcL13SIjpFOO2sYuhceYI
lGEylJ4c27tiXaw+Lh8+mEf3kra7nm+SzPTwj0Wph4Z9Wgna7BjKJCNl7N//N9dwZZgCxJgFNQ2l
MST3fTDeZ0tKD42lVtADakTZlYk2BPTkD6YIJ3u1yZYNcFUFQZyqZfBsY2NGRAlGYkrwWLI+O2Nb
K24K8t+F3ZA7P9ZsX0Fgucyd3uaNPCr7lFguNevoxuhXkV9hyoWUZ1WVwK41uTD+azjxmPcsQKyz
CP/LwsJnWVgEyDKdaPsYu97PEzbMKZkKjMGF3hUHskmsVeIr/PmGWrWKUFvYiVqTSpfiNhvwtolW
WaZpGP9oXlqWgRdboYs51mjv32/RVV9auASeF5sd2jVCnQZfibPYLrge9lKLEJISSA6bnqrfMnN9
DnkK1RKGUWbdJO9iyQAtrRoi0tgHs8Ox2LVI4HwoTKsqlSFNVXUGTEbXlO+zvjR44ULJp4rp2NyV
t7bMfCAVb0vYCwvZ3oOhcMjHxn8xO6ylea2GPsq0oqlWyrZdRtYYfn3ouhc7hRQ2tY97JIG6AyBw
H5WUuhF/sbWdJbnA3L7p9FOVxHxg9Z7j0fwWFzeg2ukj3IhvJbWBbo5+AMNn3OeXiskyLslL/YpW
Rpa/o7xof4cxAsokB5a/5YJ0htTCM7Np0zIwVOx3j588R/odeKTpKpf8E4pheaKZtM5+CSTkNOJN
7QiRfFM+CkLK4Ob9MNYkpZWNj5A61JbKZt8OoHsT3hiA6LeNTMJKocT67m87QcmgNc76R6Z00Im/
10FdTwLdV53OtQmEOq2uGjhmJFiGw9Xn7iq2X+FoDp/ymiipigOTwKMsYwnIggZyDt20zmGdgqsV
X++qv+iBwZGbKHJeYfRu+K1schuMj8Dv23t212rtBZ0YoFIscGNMxAHQNv1weDTv5Dpj1pjjwTpe
/Zvt+wRvg/LMfsomYPPYglLYxZ3PbLyemKf68QuRNglVe1pTZb+8WlmmFnKQpsPR+VYhJWc+xmGh
7fC7gGvmgMt/wn0rKqc9ZG+7PJFoUJxrY+Az52PdWYJ6g0OpSzw+MdaHWfVH9RrWM7Fmgwd/Ei0N
GT7x+OdL8EdiwAbijrGSF6GFaVZLVci4A2Y8H8+Fom9b/mcNbQe2E0vI4HPohVnhs7n2GOVkGUdz
1IQdCplYXtKags44W626NTzyYduQdxu6N3nkST9XOXIhK9cfgX63ofAepjWi7ZwDAbfxhMLEiOn+
3ZzCTbLtDDXg4t2aDwg5x/C7uGet5+knBqHyI0Cfd04YCavYw81579XpewW+HLZomhC0nS648fJ1
IBp/jiQgF3N5EcxZIZt0gajcm2t7/gCojPiVAZQUgGlrrkJYizCmB8sHSQXkOpIY7OBlz9yueNEh
fWSE2TCzTAyh+L8iZZMX4eFr40oXclX1+sdS5M7zEuws7tzVM7ggE3ZZuDF7w/e49WgYZUKUDUy9
pC+caZV6LdpAj+Vishg6UMlYMFI3wXpP0y4rLHwxNXPzYO3ghqL4GDc1PQddF7j1G1wmVEOTfRnD
QhbRztNQ39Tx3CPtFtLcDw8vn7NznpeIXeDAbZyjk2NN6nQE1+5AI2EO1YBlHRJvsZXtWLqMlvcv
VMxz4Xu11sSzesXVm3mXAePfOYnzX1jzoMdHytAtfsYuNvumeI5bkLqd05yJAlrFctJTZXtDhxsQ
MxiwTsUNhn6DUZQhvd9xCD0koP+b0GHBYqSJRVJfIE756xIEH7N+bLQuJeFTOrnkFKCPK+fyRvJk
VW1DnvTUfoBoudXUU3ifVjCgphnvm/OURNe04tYDOsIp/8R1dkxCjK4RhVJ3A2dPyzhpgqXXcjOo
iUNlsHwrzkaYvmohpzvHjgHYlNEpk7ZSDI2ouqTOM1U8pYKqT3xaNbJ10ljakZl8DmEj1uYZ0IzG
vFpax0JRjJumSaLTMCnpn3bhIrcPe3FuKaoymrMtKiAp6yRRKrcfaDKisgoXkTpbkGJd/22oAWkD
L6ZoskjmgI419H1TCHHtrJgn4wx00kRSVgMMkXsFKUUQ7RlwOfbDevUItlcBCYJGtcxeOpmD/UQY
rBhwAU26H6U2KjKKdfcuk08kMXJcOFbyg/oSypHic16CF19vmBakv7ner1waQ/qEKFg4G1kd+r/v
IEYdgBwroUThU+x90C8Zkfz27wmsACr4ghRJcHzKuIUi5fMLE3dae73tE010eVgdNawMbEzH6bOp
2B2cp2XASUJTg4BIqRNS/diBWDaMbqvTXyKcIht7RuCv1FKA92WJVLDEm6xxl0o9FGZbyy7W8iQ9
JqJjfbndLCUmEwIgF8zlWKTIuU8H67jn1W/I2i2vZJPT1nUZN85q0gckmBCH3lv+MJV1t+XQsH84
mixro+n6kDNZqnGpbVavwH3hqo/RLEcg4paUEOpzeJxPAywzYw0sf9Z+0PBNSjTNYb6FC4XnGNJu
2SUHtRMvAGqcAIKNoRp06dPRmc1dgafXxjf2tzyb8lrMR+A6PrdrmZhrZacEz0okJbJGo4CI+YHI
BAY1Yjpi7Q1TNZzA+HYhx5A5O3CejDKrN8koIyraGMusYZ6tHNsZbzUC1VQLeMv01ZhPFnMoK4sX
J2dQJgiAivov9Zo/moOCnTy/+lwdt4jTO6320ypcTvDJ8gFg+lrfXcfaFGUVJGCMqxWbH7Hi/i1h
pHnKQD/WqR7MquwMJ4+rRUAmB0ZmWvhp7VEsUocmqxqztw99BtrZ9p/7zV6P2x5U04iA+Yrm37bN
t/JO5QsNHTLt4mxwOzvng3yES/BqN1lLLeMMVzcnPRB9jqoshUtWdTWqlfx69WCIysZ6iqBwL3iY
m+HLXj318sOeZ+mad7zEU3cMbacPJ4w2W8plJjrqmXnsZHQ4oobfDwiCCdy2NxCTkQ1VwBGzJN6s
KNE1b7rm0XB3hxnj8VKAOEPdAN8gkps+RBrBDPlz8eRSsrU8nRrIbN4yvJXPV4byxouflCYhTkaJ
TCP2ybV2xibHe3vcdnFnN36EiDczlvz0Sy8OVPUrUCm0kJdSrFsXDREODWdPggjOvSX9hQHczgb9
YgXVHJHx1L0E9uPQ/VAxl+n+RK/wKJPvza/B1OtRYY48N4jJMHRfx276lN0mmdHB23V6sVyYVf/O
kqoez6Jh6AxdClbtcPGyf2/nZZUjhfeRwC1SLY8Q+FccBr/dZ0uov22uLqvnkWhwMiQtRC2Idpjb
YQLjQAdciCtuD3HHZEyIN93a8t6jXVD1FYrl/wTCUvl+2wbVwbu8pdFg+LyRHVNXQ/TjSBYFeRSs
NQ6qloOJaRU8a7otOpnayQbztJYuRPcIXfd4qalhIkFCyKm4I3Y4xivXWrQu17uXhe5VfCbygPyi
B50GJKxXi85tQ0ZM4n9EAgj+XM2qRvAA1T9xa/IWFV8HK0lXguYQZpaU1K4AaadjmqNEAyUro+Hh
C/8UBNK2qYYoEgXPaB647/7ZxyRDa9y2RVJiKx9C5acgdZyr257cbfmL2h+nJB4aa4cjoR9OhWIq
U3LklSASiMjtHpA71WJcIXR3vm9UNjKI8H3JCmYQWs9yyYz+tSdT3Ysjij50413Uv5pC95Uhkkhk
qTcDLmDX0RQWzwXf05312DnKAazCnCqBqgOKfA3CVfHPjhA+hqkeJwwWXcLyz3NWuNfbptqo6FS8
xc39DcKBKQa2UcYoDmipLkhILNYQ1xBYFzOcxGj2sAoeDoiryUjmOTaNxb2SBrnrZ/g+V20Di5lK
7qWH8jeBd1s7nouKCmZ44EEVImbnW0ywfrnAUBP7CpRT8LfKotw2mk/VncOUj69ocAncq21otx5F
NbjropjRqm8nCBoyY+70wIpiNKczubSL3Op2dtg1TLhw5p7twW3wU/GOBtqLwG/X/irbLKz8Q/yV
lZL6inmLFVddMNevbZCFyRbPucbz34ZMLLqj5B6hL6lOm/SQjvvPMvwK4tP5th39w2fPYTQCUD8a
ezd4/JKI/98KokadVTj+rhOmYVdFfrCoi3zGCVD1amL/ysZRifD+67xxtixifCs0GfpucUAK+zK3
eF16Jnvz6661dLk6cIkfZIE/Rg3aP8oQzRQI+BfehINR6uKEunm8/d1QaKAxEQ2EsNgNzjsqLVXg
1KeaC90Gus4J/Dg8CD7kZpxbmNtpw9+E67jNG7UGE8BAmQiR49DkLwcpcV8VKDQrIBcQ5sRaMgsE
rVs9oQJYgbS9j/NiTtzC1A7XwqzaY7l3ehSdRkHb0/GtDuD1oDe6MS0+mK0AybtDQL87DfZmmA4/
z1lAAZjJ1VaGjs6BTnd5Ph/4EY9DcedSHun2ntdFHBZqVjcs/6Js2WBqFFA/KP1wc6NUsAQVGi5U
/67fsFgMWGaaHnKP+Vu0IHZ6CjjCoJWB6//J1E6W51nwANVMXzHimWV6EbKI9lnVoSa9Sytr1Cnh
E7++2uBwwdSpmhH3XXL/zIZVpTj2GtMP83FgE9GlsaZxtZcmVDywdMF7jrGnQmtXft3LZf0Z3Ed4
TKBNf0snwGPy+DdnewIqnGUMDkjEFGygO3d4FrNX4Hv6mIFflJSukcq0lECXr8sv94i79YWG+Q3o
vU2xgzuWJ7DzJLVCMyP0vfm+K+ZwW3WTUXXjBU/Lzp4RtMPXvYVa8oE6XP+w8Q67vAGZIS9DIuU4
RH4Cc+UuUcCV4vhoThM=
`pragma protect end_protected

