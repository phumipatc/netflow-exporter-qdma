`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gBgjY4jdsjauEFCPquQKKR9t2H2hBjEtdHCHfEGTI1MUw/sUeI9CdHfX8bAihA/8rRrbozR/C+Lc
G+3iHEDJR8XYTpzVvR3rhve+VsWhgve6ua8JmBZpZxNJIaexF499Hu7CM4r1xwAyy9QEx/HJ1erR
HXydZOjsi82ApP21+Wi4Jf0KLK4nzOtyx9j1QDTby8B3oW8JMH4kZp5DSQ5EZP9+VU4jOoJEB/sO
F9ZSiMFbrBQEJbiArzXdkrlaMSqFwvvbdSpkAO1U7ONvTE47iCGYLc96muW07A0mF78ng3MQVWgR
0tGGjnao8yCUJIo6p4VEQMHWYebD88sDUTY/Kg==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
xg4eN+OK2tcq2oLrZyddoFkAzFEiuQAtMBfKXdAFW8pc4JailRagppBn2eFzBrVYe3hS+CBjxxMs
VY2Pe+T9JOlKbExEFaPkHQSTngsOdDBXJUyA8O5chyPFLIbci3zhJBhzIZ5zMUP+ZKMQ7DPz8ICK
1/KVLHG85wntOtlYqdJmtTcyyVtev1QivTEgNmax99TAuuxy04/DWe9y/4GVa9r33YT8K3OdkSl6
5ip0rQLszjMPP0NaOr6mGhh1KoDQgYQzCfRkRBi9JVU8ktga+09xfnC5H8UG1R+bwTk6gAdgIyIP
B647PiZgS1U33I/IjsfZEiqfo+NnVoggX5Na1gAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hMsN+Mvl2JXatY/VGxjWhBhzropOTlJq0CsGfl+M+y9o4lrNTuUN1p2rQs46M4rYX/Uk2ArSa7AV
MuNftnl1OA==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
iMXHBpLxY8YgdVFqaoxNioUtwyFCIyXA7BZkDWqdTRvNc0gE5xkDVlV5NYPlud9qSZODSUDaVIMc
RoqKzxcy1CfjC+CsUSk6jWitgPM+lfhl2JIWCr1N8ktoyZeGvFy7yuyiTV/mw//VBtWilf/Clj8p
wIFRPNHixsllqApxn/1NLqijUzOBOI0Eba8mp2js8kt97aLFUXe9/pb3HkwNlY7ExOqduXoxMJGR
u7T2TXCZtM5ex0F1e+Ktoqfd0i7iwQSeI2dLUGa7UYtl69kpO3iIMUSjVNuw74vsUbkrITwCHOXu
IpRxeQK2eUAgEaxdKRbaW0N1g1N+jiDrE8JClQ==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WKIrmG9Gs5n1nj27LEUFRHTQvp00JUCqPbe/BMzZvZBSKYvnrReoVNpd0tawd8jB4iZ9/kqDJm9s
SPDd2osCn5miPN0u90sv8VV65ugvQRiqgNOTQg3U6Q/H1t5H721ilaWSBWRBupHocfty7w/snIaE
wl5uveQ/Yl3dSGr075/F0I2X56nE1o+lLLINl4SQK7G95yw4kBduB5aAEfhuruOIKq5tjWFl3+pq
CK3p1JehTCp5odTLxJcA+D3CBPqEen++usLdxIfn6ZGEjbsU+3+qVaZZhsUNfxT9lg7VggEeeURs
utLr9cjtYmRpZ7Aejqv3YLTB0wuY6AbFaTW6MQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
EH4VK6U8XJxDZAPFHQj0V0YdfKsl4jZB7g0fFU0JFQhKY4AgI7xEy8xocPVPAQI9IlOrOJbkyEAO
qp0x1cprhvkLzVTGO7Q7JneLVhZy8GsK7tUcN7N/vur+Sp1l+U+JyjpAtmi57kvv2UqkdN6mJ1Cr
/wdyUaHu0DGoz5VPx5E=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gAtSWUGVVT0QeiD8wodvbqofQy7ivY4OwOBHu74jw1VGiYMRAlKcsY4Q2aSz7fgaUGoPkfue+sse
m3XdGXbQcWLyQjTcmH6icz9/tBSf1B0PlobFRruFbMTNtR0OOP+0y0/n6/YA33oXsrQIgWd5aifO
+ohn2S2cfiUe0Cj4ko2JTBK8kwcjBzNbLEcVBmo1yzV8mFXgxd6A966Tz6ySuoEXR7zFZsdfM66G
8EUzGTKTejLvA6es9gLXhN8KVdl+2W/8umVZBdxBzD/AXYuC/tyZ8ERmEXJKyftsUne/XGYd4eou
aD/nxtSGHshwuRbiYeF3hVfNvxxnIjbQC96Ufw==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
aSu0hIbaroyDjWb8TPL5uerF8gp2fxTR/xLh3AjrfdNAFgt2gQIfEYPiTbQeo7kwvmzLBrlC+FQu
nCNlHBi+Dez/k0wt4UDkEQT58ci9fUgVUxfoP1bs44WgP4J5zBpavVoMRDCYBt0dUmc02mTKR0vD
XkuxxWIuLEP7RiF5TMN9nzXaOv8suoPYTzUlcHEX0nOMLk6KsCXekiQq7XVLnUb852yw1iMQEFSD
5oXn1itxgaNoRh6i96roHlWjkPv2S0BzBpL1Axl6ZPjCNuzOrYuvh0oGoSxDpgNBYv790d4QsMT2
Q+hEX8vblA/jsGsG5hWEFsS9bUyvhsJZYZ3Z2g==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
pcyKZrCeVVyT8hJ8yXv25ithF0nCG7HTulBO8t3ZC+vU4KaHJqwnagwqDHBugxfOy1wuce+HJptz
eBijfb8MbvjNqOPkgvhB4WvZgzyjOxaCBV5EMKng9KDEWaFAIwrPtDo9lvCn2Y7HhrUw1+/NOgXA
pZiyVVxTkbbzrEIRt5I=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5j1h/tzviXGJwQm71UvYLal4V7trnhlxHzbA9A+Jh0reXqaSLSBvNai468zw+r5lMcy3wFYxIMK
c6on6AmM0cAowoI6L9/TLu9p1i45xkpxaiE9VtQXf02BvzL1YPIVFTI7i5F7T4XimtlD3ejucnP7
iJtYUsLi3kDkyy4+R5zciPg4Bl1uG7K49t5TkD5iUxhxbP1Eu6Dy04WQFt5k+bHxxYIPPooFRJzx
yEKPJ9WQOY5rdVQt9rczjw/zEW4pMFGMBICnaJdWvD2lDQpClV90YMfEUuO/zQgqulh8gNS6/Vgw
ijWhHXbxTZ3Oc1TCuWfrwSTAaE2nW9/1QimYow==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2912)
`pragma protect data_block
ddRdsf0OVem++Ihid0l0y6R36MxRFUTWwp/1CAdii07rSAprP46m8jkiGjsc/804/g7VgCsvxTIh
imBuUABCHJC25uWE08LOdDj7VUk10hzX2UXCNEcV41ENSoXjlz+Oz7gp7as5+hUCetp2t7xS39op
2zInf7EXpGoTZa6RjVlFplM/0Vk9cCBh9RF9vTWq5imGBZoftE/ybucia/Rj2FvVHcIoeD8mpR3r
0zB5o4eXpC/E3102I+sw1pxgATzgDAtBqAtBByGrT1sk2FJL1D206DR5ORZ8bPDzzXoh6t9pFrKT
DA3BnU9WMg59YrfxPJQsQ7TyCGxWUWj4jph3s5fRW5bnYcWdbKd0lJkpapr0vhtZZAfHy+iybPoS
OpWorcVtMoj0DS6tsxl6NJXWuShXtLIrpHaG395uHHWkPwoW+RhqLFyDROKk3JOtcUbpHFG6O2nZ
dk792OhHAcy8f9xNWWMs3xRB4iYe+/Dn8mxcbbaTJa9xpP5y/Pp1+qfZFnzpFxXoVCz+OR3gO+SL
dNpj2u73d4tGx5dsywBFX7LrXF87bNISJIPbpbGVa/6f6A83X7FaydzSQlEGjogjeNteLcPcayfq
zrjfPNLerX5Y36/QdM5YKbOaJYlf7NJtDpHft5pLUj4phQmj9ulTuXzVduf3K87bqCKU1h6Z67jJ
pasSI1Hh+U6QPwheqwzy9Y0DtW+Xs1c2Q+jCmhIlq8IYhLK8jLA8/VaEJdnOEOnfv2lyc5HMI18K
UfiRhSlOSMeQlKYXzpn0jWd5ujc5FBG3kxKxhK1Csd+vKftVoGzf95N/W3NSUmqcTendaWY3nzwW
yPr/uRN50CO+l6D+FRNcLhV0zw143pwQnvBdnzd5Q9n+HitSZ14yJb/GNP/kwN3HPVvVF1NBYWJR
7BxiJK+95MOm/SUMt9MEX0g9BA2wOgk/WWXJdr2FjRlhVaIzs5P4h8Q5nn49WXT6+i5en/2JjyKi
pa9D12j2HKd4Y8nR2dR7ZmbTAGmRucfJZqlSrxCNuq4s/bhKO6XshaeFYO+u63M+YThgMgh2EVS+
BtWYzOO3ah+n4lRo0kB0e9TqaNsLqnf1YLyKYEheBgBxD6s+CeHEkCeTiij5fF2cPZcKxt0Bzwva
t5q/Ssj+C2GCWUXWaPExZlxx5EEwC+UZm7LAgI6RCMp0AAQJCgSnBEhP8F5UKT0fFl4lhH66eQDu
Is3u8NpJSwpGuuMcB65kJ/DApW4prTUhGmTPsS5inFZT+/neyY+CvjZ3WS15tZsWRFuciwmemT8v
XvagXxB7Qn8+oM4abCHR0/RY7VRaP3D4gsi+mo1sYjGaWrYjNnXvv/D2q+YVo+TIbONPb5iC7oZf
UDFgpd4v3oOr+BWXn1ogHQxQMzg4E/xiWmJcXdJsAosyBUP2BO18SaV7lI/tARAJzhhXJ8wPw1TZ
yrH6UpwRjSV0dDnnRWjnDIEP2faxV4G1ApJNW1kfMnzlIo9UhJK/j4KsZITo9z4JeTAWVG7GTvyF
Ml3o03hRqsxunjxc/NS3sAzpx4lmB9KyhKKTN4hdVdHsVzQei06qhDqOAMvS4LiTAJV8x99dMUzE
X0YCu38hGE5qEY3jcSBidCuOb5BsYDZFuodFLgBUdCQ69c1fzJmo6ErIPGOnOiTssz9KBZuIV9dI
k33MIUaAe5MTZ8fRooYFxmCUPY60yFon0xVd4N4syiD1U3RGomd0UfTIFoPfLmu9C17eFyEpH8ZK
hJ1Zw4Cx0detVk0ecs3ECyBvLewMQRMiTJAHZGdvrJLUXnQddxj2xgtXk/WTDJ//khscnuOG3QvH
rHVOsR08tveoXwyzV51slIv/l2ro3+OQGLaMUx7+rRE+84CMDSied6lHVH7DpifVfPoAsU+UR+E/
HQCR30TgNqlzdMHJehPGf4LOt5AF0UB9CV6XFBo65iJEmKBVFb4GVL6ORaGQahCkl3AMjPAuDWRq
8ADIdfQOGXZCzLtuLRGjqaiWEvw+z59krI/mhcJ0K1Z+5aOh4i45hMb717EFtOQAMzLPlvnFEpPl
oYAzgm2bpxy/jTY477SZ7l5ZyZDmlYC+oJBMexPwGAK3tozF0x4beuGKseRdPYBdDL7VtgFcpZs0
/2sX+cgbjm0Zjl90S9SIHEHk2n/3aBsWcC+cc3yakB8Sj6ATFHuzrF+GrFX/xGYOczw5vMWarTvS
cYK3UpMPYvm7m2QzkULu5my6ZKEX6Cve3ev22vtdeFk+SL/rF5s9JIboiGKZQc5DHaczexrSbziY
nQpEjGaEq+lcjpA7QOYTK2YvrIbiM2RmS2uhWXzmJScgsc1BVPjeWraW+B8hQJAcBEYBNqCpZblZ
CfcJn+QXlc88l9Ik5qBItvS/N8TT3DFPAv8dOdNrccJMEdEENV7lyu9y0lS5i3lXxV8V/+U8tBSI
RSa9LIGGTluJOYf88xJWwBKMU8p1k1E7FNLC8ZZFMwk/PBvdS+BiWRnxpmBMJk1MgkLCCudnC4IZ
claoHCvo6wFyKcbewrldTPupumAT5wbruSb6hGFEMm8f0wwmF8fZGlcc38ayT14OcjKOE2ZXQ7hY
L98ZaJWlvtGkAEwvBpvKXXR6TJCdNAXLxmh3945zix5y7eB2M/TT69ZukORqMBVbL0vDw5JsCkfH
NFIbOo9uU/DMkgGEehlqEkZoE0diDSbwx0k3h1nY9MYbPC08vkHzBWkPs7gJF4EeaoP4t9ehTKA+
M7tMnhUvgTzVNR1fDIRonZA6kMA3Puuj6YVcX9Zkp9dORGCkcJVpUI54CuMqxqiNwflVdhxo56ew
qsYWv5uaS+X9OIwAH1a8wXbC2aDrPX/s2eVkbB8flHMRdctEzmJqIJfNNoz+lXCuV7G98z3cQG32
NcQyF2qrtkioGMzdzqShWgZ23BbPpuXdU8qux2xSCtaIO9lUIsqa/zgGeXoBaiT/m1dkYMSz2T75
jwL6GeWKk5YKzFtBWFZHX8dXTorvL5d8JsRqJIUrpaRUVbKxCySlvPQGDpa8hKe8fMnpMWZgWxZS
iPbnj25i29PaT5VzghhbIIhLHFkyj3vri3dnCLKdM3xMPfAOFPN7iaGojZzWz82zzkBqZ/ICBqBG
crCNZYsJpFKnpi2akJ1cV+C6Sn0zj+5JFcMp10pT7nj02zRmKEOT6lNRufEjB48BU9KQqisZKcx2
szhX3xRXV0/ULh6qS1VHIkGxJsNyn31GbMkoVjpQ+AbIc8tQJVdiISxrulDp4Od5sP4qFFKunGFZ
/QMXGu5J4ZfjIy+5Fb0lk14gn6JAouCu0kPDWCfAOzdv166HzjNDfb0DtmEzZEu+CcwQs8qxwsP/
/4KuH3nXqNyFfp40vgGGGaS41aR1XOePAZxYpFAFwXVqHYJ1hWGP9FrrgBJlYm7lSJP48+8a99OQ
lDz8if7NEPCC6u1JXJofYcv2tZ1MFyoTY8Trqt6/PvwFsXm9jw6jTlTYBm1p97aQUcJurXVbvq9s
sLqp/DWBxAfxpNsxbGoe8QikvwqH+IVPLxvtytBmlwDds6ouMX+TyC7I5SPEMxV84V9Xb/1dKFtm
Mc4faqcISCxXOisCKKDYzAGAaJajJ0aFyop9gVQ8oqGZzq54bxW/g2S7MjLwcR4tLaAWluiX4Dnj
1Wd9ur2wlJcbNixr5CTvcMG4oAezLIL6tPZNnTA5DwJPzr8NTEfnK+K4BHQL+p7dGnaKEzuPWcbV
mJLWcPTt0F2hiQxbYCFSXi6NZtWlQweeNalJQ6b6y87R5vupjfchZ6Hw1eHgQRBggpsA5V8Wb7GF
T5WsjihWvJmeTHh8MGIJ5ehZIXDRAKU3L7OoMGcnA4fXpUUBYXB7bekaAYngJa6EZlWbAKZpzTEQ
nZdM/ss=
`pragma protect end_protected

