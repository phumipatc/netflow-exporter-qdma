`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jlgGOAB9z4WRhgG27PxzR2C/U0zMrA3PmuoTGKCjWCt407sXMKGoGxrQdP1pHGBMQMj5RV+pzC/U
XXK/Z2kiEzbGgCkB0XbUv4RkS/GJFaC/2Jq/C1KDFUJZThKe0a4oWZoAFcwi22tXp6GXrss6QxGd
r5S2mAEDe6WDlThYvPuedTpbKZfMWRld2oBweLBdGgBqv9QrYVDGHliPFHFmYn94TVcWAeoC8aGT
NMuPAut5PDeWihTt0fmOzn/kX0Zb/pCX+esj7B8W+CJjfSVnx3gtB9HoAfXSwAc5MAo4/Y7cFaZV
UMlFu+1mxfZGpECx3gN/BQwiUwBis1NKd1wHdA==
`pragma protect key_keyowner = "Atrenta", key_keyname= "ATR-SG-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 384)
`pragma protect key_block
pgoIurua+UA/tTh8OyCDrs0t4Tqn+M7A0WTUZomViyshGPiGTzfs/9wbWgtkozEPbtALy0Opnt5p
Ah+7I84j5aWUHZ1nxeE2H111AClC8mOw+GeThxSH553Bym4tcl1HH39WTxNqXaEN2qecI7T3DSXu
Kc48qubYkcy700drbjKCVB0a1SPphnOeHvKQ4bdf9EByYGew0Huw/qsH5t5dEPPLIDofmyIxwKpz
zBxZYQklV4tlKQPCPZqLJFPTKsjEUQIE+LxsCRltPTAdAxk9gQtBPtNAKOcEYz/pBngmHiU6w73V
yX1rutLwYC4sT7dIHToh14JrmYAtbSQrwztGngAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
gPKH6w1Ih9cmSLsX0U2vvQHwExM3dZEZZ2fO3abwkBRKFcIkdemZm3YtlJn96I5WgKHYdhUPwMZ1
9irO4O5T3Q==
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "CDS_RSA_KEY_VER_1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
JVe8iqXaJQSF+27lIaQTQYDIJqRIUDpaN0F23c7BxGL4LoL/0z80lPb0d179fV/RXo8splRaLPSL
4kMAXFsF7Szdxu2uwvuON7mP2Z+b+Wr8/NY5U/sy/o2NA+OULVRbSWUPc428+UXCmJP/nL5cKMoy
mA8BBePbzFL2vhqUq5gJsvlAUziP3x9xiMF8YWkDnruJYwXHp0RRomEpuViMU/vDUfFGMrq8+Ukk
ubGKzUyKD8hIzlYtIXo/B4P43k0Vn/b3tzqI2EzJDX1o+lAnTajLSjEvzvknZJ3/1MYoZjqCcc/G
FmsArhCXi8FUwOYmRTtZoGoq7jICEQoV57582A==
`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
dRh0wEpe9Q7ywStO6dM3GOdF46mP4B6vsrLDK/5qys+sHftGU4qmN0bEZ/l9y+Xjh5+MndIzY/Cx
z2TcdnQJXVJxvb9aK1E7j05cD6iI5EYExEHRjQv6e1A1diESh0S68HTz/Sb4m5WedXIfCtD24wYQ
vmFBUBuxWmTLsZSAzR3+MnuClv3t/H0igQx03wdvrOqo6MRkxvlEoE1ABJdF/Jt5V3vo+ZQRQZ3t
Qq3b2BrzFcTP1gQ47EzvQ3n134JXDg/QrVp20QAhBymxnVEjmxGxIjjYK+ruPZpEvy31nH5N85Rk
Dva1FIAH9nrS5dunfKYHWrKKlJc3Oh06rTtFyQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
uJgByocPfRLHu1Y3QyMCqx8S/ndi0YZN5UbbuosWLxEuh6z7maiuCuKHILU4PHNdXqbq4M0GysE4
27uEQCP0Isib/SUiwuCL8qx2By9ZWWbBTo1voePp+C+M3wfNFDzARKfJOHS1coM/UaBd7TMLNYiY
vgocVI7LGmGgThNTMXM=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ekso/C6zfUdLMQ91OSQ5d1MUIDzEwd6eWoEvkhZ24GoU6P5OoHqboGQCOBJqyEAAHUfI3nM82lFy
s96eqFNewSTVvrbaXRfiE4X1MrvQS5oRX2jQc43Y7OS/JBhdXQH7mXJHJ/UEM16JxtDuTdvOoclZ
RBWkskCkfRWXZyz0PCRkFz1Gu9Xr9v0JJCaFd5dkTZb8Jfymf44GdXWJ7Vl8t2C13XSyp6kjr4+U
KfTuYkDh6dJmHLbsjDJ3p0NovNeld9m0gbAL6RUBmP5fWkMPxhoajlH9I9cf7l0BU7HYvepzi9/d
gSRGTW/nyNtDe+mySfUt6QHf7jHevdDz5mm2kA==
`pragma protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
k+afSPQkIbMZ6jZD28uTRocmrVR9Cas+g94EaIidrLGvQgTgH8aAd8WD8H3fNDcCvGTdiIBMxJST
uB5vcZXhjoMKNYFVmaJ7oFcJI0NcBjYSc07Ark8JCjB+gNS6c5mBEcaTStiDe3+E6OrJcRbafqlw
WATmDDrvgn3Z2b6FuPUdAXt1Mff9ycADUSrXuerZOq2gYVYeNrgVF9ze/+O2cy/rb7dmJg4y8YwX
UGNNxowL//zaM8DKDkBpDzr74FqNHOE2ynt0OdkyZ3yQsFSL31yjNpVc3nwA+gnNLaFDhvQLI54p
evCL2rJpZritkMMwrEMFgNUVr93///ybDb/Pgw==
`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XB/bUIV8R/4buqyO0MxmNC/moo7OikXylFfep0rWRgHgdzKqXX0t5OoEg6gqqb7M+tHlJhfVAFhR
YluDe1Ixp6Tp3rkgfXgY1fK/R4sjj/KDyBecn33cZYOWEwwh20RcjHqtZmzRPPJP21FKmujex4lL
gw4/+PUk1cjSbmTpX2U=
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2022_10", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
oldieGkvKb9DASBFBVtk3BR1HO7Skcj6QrqoR8cONL3Jg9i3GPl4kNfPS4Dhg+K2rCVaJ11/ulP6
Qkb/nDvg9bxwxdJHlCk2k0WUjtLyKDeDpLpOKA1Rgg83XpFX1NwIuZEQAN4tfIUANfX4/gaHBJm6
LJ4+17PP6MUs3wxnwACfxHDrxYeOXqBDzoC73uTfZxgnBy3EY522mrEmZWVQffjHRLJLkdBtBZRi
HZXVclLxBJJNqTBVJkhBfR69kaIvmnjz2/tJCAYcuOfHHg/mvsMyJTv6otJnVTbSZgkiQAYpfbBR
CAUt7zlvO33pD6SY9H0sznkRzJUUDXzNCMLvKg==
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2912)
`pragma protect data_block
0/CQP4xLIwggsxczTWb1d0wGItQZEfDbXvhwpc3Qs8V/2tdaXL7v9MuCSR3A2VaYqwrsJnlUGY35
aosFHfPF86/UQwd8Ce1/kuWKqGQ3qMF6TEIAviOY5i0v4EiyCKcDyyVVEoxz3zsWeWeaHWMVCCuM
uVpAuOJ0Au+VjxFXEX5wMvHCem4pKfztYLc3h0qCaENLk9JmfvNzaMRUpDdGN47MyAjmCyN1tXMb
B0JC5ZUrMN2yOy5++PS5tfWSfbVXH5ItOckYO+sisMvRk37mroLt5eLNjkBGI1t2m7wK8w9i0Fn0
IrVpJMWrIZO4EQP3f+vXWgvJHFBS5Xq0OxZMcXOnj6RuDWbsL75BSTeuQ+PETdT9uX2piIG+6WoC
vUtZzQHJh+kJ2PEto8nMVx74EeNfThWggHpL4218Qa0lB9ktlRzrMs/i8uD03/f0qogTIVFu+OVh
qjudcy1d9HtZLmv/nWCbuFpipUk4Fom6aG38zk34Bv0Q6R5A7/CHo09eTtikgn1V4OswkpTtVt+J
01ER8BE3Q8aeMwaJaC75rOqwo3JFQqopOMM9tPudb05ai3HFtZKUYnP+1HUzCoLIBtR8G4Ldsha4
hmZnHZkemOen/ra69YHLjgjq23AU4XwbHlopgPD3PPBHu1v6B4kci3m8l58hO2h22c+RKMXxb9Zr
dpqXMVVZXtSojCmKNHLReAV/RUz5WfNZBNY3Q4FZee5M77smH+GElQw7j3L8hd5iK6wkRyxKE+vi
mwvufQ1E6P0eXFvElME/JO4dfXDyXfeRi29S6EMD8LOSx94eCXbV+08z2clFczyA8iVh2CY0O8uf
OeTvBP28SAk10CgiEKHZve/hM7LUigHQqfoqkaajyzIQFhJ2hmf+EUUUpQDyflgZ9gsB1zuTjtH9
b4mKR15RXUtFt2Nw+oZT6Fjm22VesqRP5oHc1fQT3lbXbAZQO4oExAA9k87eQxXtUlIK2ktIfS/a
MOGjwfpRTgxr0GDIPXtA1Kvt5gg7Ct/18VrkuTe2GWx0/lJ4WYELbTTUzRaFL/ECB9qfH5Ev6p3y
H+2gNSov/xiTkuuAtinICHbAz8W8ML+TFCE6I5FSWUyH6ACqHaRhs6kuEP76Ddug+vOTIpYLJSmY
9owrtr9RZsro70eFwWBLMSH/9G6Jk5rBamjJusBIqMaLrCj54eNV6hWP86oqntnet6V+LS/oSHS5
5cXvWYwZhO834tdrs61OIKq/Y9H4XDXXj2/cJUTMhH3SSquyknOCOC9chsf1Xi6EhlpFUMDYLErr
6fEfGhb5wiawL23GvQaI6em1f9nkvKb0mUGf2L9927qOTiJxWhAFrNakcsIBDGxq0448w59rLIUX
QymKhl3z2uEHjvZhZnaQfGZXSdIm1IwjfRaT2XdXcb0VIIKeXTMyTIz2hh6Qhki1Ppt/dp0rR4DB
dYecr+fXSl9wUUCDtKflrKIuk7aZOCvFL7Z1l7F1k1wB+i2dcYy9tvvd4c026UKBMSN0C5b1BPgj
zaOSe4djG+iduqgIZruYekVJdwZbq6Ho1cN4BFA6B3DjTtgdJBLJCTOCqNOFDbvOLoNqv3PdNV+l
DvQwoKHPIrl4jGeRjyKL1wYZIThv2FwmyVkSKb/FuClRt+ptIAVjxMk4iG4tqW6p1wEs6rT97p8L
Zilfm16SClzQLeTWfVtoSAF+XTclx2LvPg7mG7tY5dSgA3X30tRb1nk+e4qQFJihaV+KJ26Lazvt
EbK2c7LY7wyWjrLL+8yqjYVcpJdEJ0D7c26Fd4OlD8h9c++A0+qhs5PxPdd2BNXd38wGoTQwHcEi
1fREbVd7PUSqQpafrRAQsrhLZbopt0/8UZYEpLZwt6YvPDltxQcXkwVQRjnI4ajRwel4ZzkGs/kA
cS8gV06yujeATbFovhIcUXVLUJ5ulQUpYUAFCjeYlPFruhadXP8ia72o4xkUSgfJaqZm80mBEjeV
2msEMMyvscCaEvX32WSuqCkAEMG553m8tGmD/sRX589fIoASWYt6TmzFMSebTPw46qdU7SVx+1KE
aoBhgLClMx9CyUYkOafSbIywMKaToGetFbFCUM97paidCjWmIsQj0+ykoJ39mxNUnCbbcFIzvJy6
nErvt5ebVMl9/c/04GsdxTDl75JpDz0cIsjOUUo9G8FzPQdLJYpdlSnwk2zfzm+SIm0vUkB5O7qM
VjfqZiuPMjdHw8ggJbNy0v6JunYwBKiVB+v98RZPOipKw6wya2fQ/c4nPWCGrB9uEHrURv0RpOeZ
XQJi37xUeXMtKc4VjE+lj0Ccj04c7VLONTepA8D73jcIzr+2jRJXY5SulHyc30ASlWuBNwRTMxjS
3VZgkacrm3NHXty5XSmKiBsLD22dbmXjUAo5hmjicMbLlcF0xdxyF//QpUuDNhcVl/b9lO4sH3L0
Ub8LXRgfidjgvQdmgrvkmia8yGgoss9Rbnk0bwEmlRrXAeRtbmVsLny3Q6PrrsI4L0qKCAzNT+Er
TvBv74y9CGSoFKoVipaFAwqD526uJ9GCFzLD6lFVi8tx2SDlyxII3RskRKmi9mdaS56+EgZsg+0G
u6fTKjXW6zQS1C4515a7HpfwtwpZdKdBl6eD9TVKKSpcpyUVfAtEQnL2t5nFVi9rurSDDPj4e+VU
qYuN0rIfpRSUwgaaaR/+qSmi4G9Xeg0gqZVCxVu9GMdrARW0qANz2c2J9j5w+s/3ZX6b/OBYn0Qk
4KKlHgM035ODutDMpR+yT+7Pud1lGxDU6vmaTrp6H1Q3lE0iss1GMYPRht6+/N0JcHUYuBbqCqnr
pV6WduX8FDapJde1XQUuNXwow55DgOj5h54i4gE6nF5Y86R7dlRMe6EDrzfVPoDac6S2+o2hHSrg
+NgHh68/2Q0AaKdatjwxM9bBqo3LXxXcz1YojyhXryJJFeb/UlLzly4FIXSUzWsV3xZ+UnKzs58k
k1h2b7CN2npZhwBObEGjPDZVOFbQEC/VECwYKLctIig0TBNg0jNsayG2mNvs3XGtTuf28s49s59j
OUaatbUzvTlET/004teJMMl02V1fllMsXAPO282i2fNS8xDHn6KKwcF/18sQq5PRiuXOOI5XfIy9
I/jfZVsD3W+MooNIn+odce2CUfk50M2AsQaI+AlKnjMafZn8WDNSepFkbZD3XrMt5R4NbI1gzu98
1cViAkgGApKUxyFXn5a886OgPl3D4eI4UFcL3S1vdFufUREBY25VcnYqNVr8bUpfG31VQw8d/aOK
atKhU7gzqNsdrvrN6n689NGuibXeeeavd1WJqH+U0Snth6xvDGOAFgGo+A1YOEZsI/VSuVGjxe7r
Kxm2AOvGGFV4EGg5mebHXzXZdfm5Q0bdSWtcevixqWTmoHZ/1oBxPvEGtAyvVb4JLFUlSEh7blNj
SoPkTp0TbgMfmRue23xv9J7Lab3Isp1OacMiRHAhhg8w0H8S3SUA9pgvn6my/h9IXOiBDt+bCgBU
sZmzkt8pXwWGGTIZ/nRaf2yFSI0RKj03z4fYrRDe4C9rIu46na5IH+AjDwNu3tThX4qv/nmsJ6C5
DOPt/+6iAS4CXyBX2s2LAsvAShcE8izDRBDJ+SMOLgxQKFvoliFQ1gZ8FqwtNX1qGse3ac9EFf5S
X9USuW7WVkEwN50UyC/bB0xo131empXYDPT3UMUdDvLCStOrGz1L/a4TjspSsFlqzeH2D1dakxf+
bEWCzsSSE1WmH1o8+yi+3wCUxCUgRamANA2CnkE8TXwwvP7z3l1Gl1urYONKIPeO58ku5vJAFsmK
HNjSI6EEx6DOLByH/fmQaWoxaWSujyw//8EwnABNEottYWM50AjarGr2Xx4gQ0s9JiB9ItMEwozf
7U39Fr8=
`pragma protect end_protected

